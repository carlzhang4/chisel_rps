`timescale 1ns / 1ps

module tb_HBMCompress(

    );

reg                 clock                         =0;
reg                 reset                         =0;
reg                 io_axi_0_aw_ready             =0;
wire                io_axi_0_aw_valid             ;
wire      [32:0]    io_axi_0_aw_bits_addr         ;
wire      [1:0]     io_axi_0_aw_bits_burst        ;
wire      [3:0]     io_axi_0_aw_bits_cache        ;
wire      [5:0]     io_axi_0_aw_bits_id           ;
wire      [3:0]     io_axi_0_aw_bits_len          ;
wire                io_axi_0_aw_bits_lock         ;
wire      [2:0]     io_axi_0_aw_bits_prot         ;
wire      [3:0]     io_axi_0_aw_bits_qos          ;
wire      [3:0]     io_axi_0_aw_bits_region       ;
wire      [2:0]     io_axi_0_aw_bits_size         ;
reg                 io_axi_0_ar_ready             =0;
wire                io_axi_0_ar_valid             ;
wire      [32:0]    io_axi_0_ar_bits_addr         ;
wire      [1:0]     io_axi_0_ar_bits_burst        ;
wire      [3:0]     io_axi_0_ar_bits_cache        ;
wire      [5:0]     io_axi_0_ar_bits_id           ;
wire      [3:0]     io_axi_0_ar_bits_len          ;
wire                io_axi_0_ar_bits_lock         ;
wire      [2:0]     io_axi_0_ar_bits_prot         ;
wire      [3:0]     io_axi_0_ar_bits_qos          ;
wire      [3:0]     io_axi_0_ar_bits_region       ;
wire      [2:0]     io_axi_0_ar_bits_size         ;
reg                 io_axi_0_w_ready              =0;
wire                io_axi_0_w_valid              ;
wire      [255:0]   io_axi_0_w_bits_data          ;
wire                io_axi_0_w_bits_last          ;
wire      [31:0]    io_axi_0_w_bits_strb          ;
wire                io_axi_0_r_ready              ;
reg                 io_axi_0_r_valid              =0;
reg       [255:0]   io_axi_0_r_bits_data          =0;
reg                 io_axi_0_r_bits_last          =0;
reg       [1:0]     io_axi_0_r_bits_resp          =0;
reg       [5:0]     io_axi_0_r_bits_id            =0;
wire                io_axi_0_b_ready              ;
reg                 io_axi_0_b_valid              =0;
reg       [5:0]     io_axi_0_b_bits_id            =0;
reg       [1:0]     io_axi_0_b_bits_resp          =0;
reg                 io_axi_1_aw_ready             =0;
wire                io_axi_1_aw_valid             ;
wire      [32:0]    io_axi_1_aw_bits_addr         ;
wire      [1:0]     io_axi_1_aw_bits_burst        ;
wire      [3:0]     io_axi_1_aw_bits_cache        ;
wire      [5:0]     io_axi_1_aw_bits_id           ;
wire      [3:0]     io_axi_1_aw_bits_len          ;
wire                io_axi_1_aw_bits_lock         ;
wire      [2:0]     io_axi_1_aw_bits_prot         ;
wire      [3:0]     io_axi_1_aw_bits_qos          ;
wire      [3:0]     io_axi_1_aw_bits_region       ;
wire      [2:0]     io_axi_1_aw_bits_size         ;
reg                 io_axi_1_ar_ready             =0;
wire                io_axi_1_ar_valid             ;
wire      [32:0]    io_axi_1_ar_bits_addr         ;
wire      [1:0]     io_axi_1_ar_bits_burst        ;
wire      [3:0]     io_axi_1_ar_bits_cache        ;
wire      [5:0]     io_axi_1_ar_bits_id           ;
wire      [3:0]     io_axi_1_ar_bits_len          ;
wire                io_axi_1_ar_bits_lock         ;
wire      [2:0]     io_axi_1_ar_bits_prot         ;
wire      [3:0]     io_axi_1_ar_bits_qos          ;
wire      [3:0]     io_axi_1_ar_bits_region       ;
wire      [2:0]     io_axi_1_ar_bits_size         ;
reg                 io_axi_1_w_ready              =0;
wire                io_axi_1_w_valid              ;
wire      [255:0]   io_axi_1_w_bits_data          ;
wire                io_axi_1_w_bits_last          ;
wire      [31:0]    io_axi_1_w_bits_strb          ;
wire                io_axi_1_r_ready              ;
reg                 io_axi_1_r_valid              =0;
reg       [255:0]   io_axi_1_r_bits_data          =0;
reg                 io_axi_1_r_bits_last          =0;
reg       [1:0]     io_axi_1_r_bits_resp          =0;
reg       [5:0]     io_axi_1_r_bits_id            =0;
wire                io_axi_1_b_ready              ;
reg                 io_axi_1_b_valid              =0;
reg       [5:0]     io_axi_1_b_bits_id            =0;
reg       [1:0]     io_axi_1_b_bits_resp          =0;
reg                 io_axi_2_aw_ready             =0;
wire                io_axi_2_aw_valid             ;
wire      [32:0]    io_axi_2_aw_bits_addr         ;
wire      [1:0]     io_axi_2_aw_bits_burst        ;
wire      [3:0]     io_axi_2_aw_bits_cache        ;
wire      [5:0]     io_axi_2_aw_bits_id           ;
wire      [3:0]     io_axi_2_aw_bits_len          ;
wire                io_axi_2_aw_bits_lock         ;
wire      [2:0]     io_axi_2_aw_bits_prot         ;
wire      [3:0]     io_axi_2_aw_bits_qos          ;
wire      [3:0]     io_axi_2_aw_bits_region       ;
wire      [2:0]     io_axi_2_aw_bits_size         ;
reg                 io_axi_2_ar_ready             =0;
wire                io_axi_2_ar_valid             ;
wire      [32:0]    io_axi_2_ar_bits_addr         ;
wire      [1:0]     io_axi_2_ar_bits_burst        ;
wire      [3:0]     io_axi_2_ar_bits_cache        ;
wire      [5:0]     io_axi_2_ar_bits_id           ;
wire      [3:0]     io_axi_2_ar_bits_len          ;
wire                io_axi_2_ar_bits_lock         ;
wire      [2:0]     io_axi_2_ar_bits_prot         ;
wire      [3:0]     io_axi_2_ar_bits_qos          ;
wire      [3:0]     io_axi_2_ar_bits_region       ;
wire      [2:0]     io_axi_2_ar_bits_size         ;
reg                 io_axi_2_w_ready              =0;
wire                io_axi_2_w_valid              ;
wire      [255:0]   io_axi_2_w_bits_data          ;
wire                io_axi_2_w_bits_last          ;
wire      [31:0]    io_axi_2_w_bits_strb          ;
wire                io_axi_2_r_ready              ;
reg                 io_axi_2_r_valid              =0;
reg       [255:0]   io_axi_2_r_bits_data          =0;
reg                 io_axi_2_r_bits_last          =0;
reg       [1:0]     io_axi_2_r_bits_resp          =0;
reg       [5:0]     io_axi_2_r_bits_id            =0;
wire                io_axi_2_b_ready              ;
reg                 io_axi_2_b_valid              =0;
reg       [5:0]     io_axi_2_b_bits_id            =0;
reg       [1:0]     io_axi_2_b_bits_resp          =0;
reg                 io_axi_3_aw_ready             =0;
wire                io_axi_3_aw_valid             ;
wire      [32:0]    io_axi_3_aw_bits_addr         ;
wire      [1:0]     io_axi_3_aw_bits_burst        ;
wire      [3:0]     io_axi_3_aw_bits_cache        ;
wire      [5:0]     io_axi_3_aw_bits_id           ;
wire      [3:0]     io_axi_3_aw_bits_len          ;
wire                io_axi_3_aw_bits_lock         ;
wire      [2:0]     io_axi_3_aw_bits_prot         ;
wire      [3:0]     io_axi_3_aw_bits_qos          ;
wire      [3:0]     io_axi_3_aw_bits_region       ;
wire      [2:0]     io_axi_3_aw_bits_size         ;
reg                 io_axi_3_ar_ready             =0;
wire                io_axi_3_ar_valid             ;
wire      [32:0]    io_axi_3_ar_bits_addr         ;
wire      [1:0]     io_axi_3_ar_bits_burst        ;
wire      [3:0]     io_axi_3_ar_bits_cache        ;
wire      [5:0]     io_axi_3_ar_bits_id           ;
wire      [3:0]     io_axi_3_ar_bits_len          ;
wire                io_axi_3_ar_bits_lock         ;
wire      [2:0]     io_axi_3_ar_bits_prot         ;
wire      [3:0]     io_axi_3_ar_bits_qos          ;
wire      [3:0]     io_axi_3_ar_bits_region       ;
wire      [2:0]     io_axi_3_ar_bits_size         ;
reg                 io_axi_3_w_ready              =0;
wire                io_axi_3_w_valid              ;
wire      [255:0]   io_axi_3_w_bits_data          ;
wire                io_axi_3_w_bits_last          ;
wire      [31:0]    io_axi_3_w_bits_strb          ;
wire                io_axi_3_r_ready              ;
reg                 io_axi_3_r_valid              =0;
reg       [255:0]   io_axi_3_r_bits_data          =0;
reg                 io_axi_3_r_bits_last          =0;
reg       [1:0]     io_axi_3_r_bits_resp          =0;
reg       [5:0]     io_axi_3_r_bits_id            =0;
wire                io_axi_3_b_ready              ;
reg                 io_axi_3_b_valid              =0;
reg       [5:0]     io_axi_3_b_bits_id            =0;
reg       [1:0]     io_axi_3_b_bits_resp          =0;
reg                 io_axi_4_aw_ready             =0;
wire                io_axi_4_aw_valid             ;
wire      [32:0]    io_axi_4_aw_bits_addr         ;
wire      [1:0]     io_axi_4_aw_bits_burst        ;
wire      [3:0]     io_axi_4_aw_bits_cache        ;
wire      [5:0]     io_axi_4_aw_bits_id           ;
wire      [3:0]     io_axi_4_aw_bits_len          ;
wire                io_axi_4_aw_bits_lock         ;
wire      [2:0]     io_axi_4_aw_bits_prot         ;
wire      [3:0]     io_axi_4_aw_bits_qos          ;
wire      [3:0]     io_axi_4_aw_bits_region       ;
wire      [2:0]     io_axi_4_aw_bits_size         ;
reg                 io_axi_4_ar_ready             =0;
wire                io_axi_4_ar_valid             ;
wire      [32:0]    io_axi_4_ar_bits_addr         ;
wire      [1:0]     io_axi_4_ar_bits_burst        ;
wire      [3:0]     io_axi_4_ar_bits_cache        ;
wire      [5:0]     io_axi_4_ar_bits_id           ;
wire      [3:0]     io_axi_4_ar_bits_len          ;
wire                io_axi_4_ar_bits_lock         ;
wire      [2:0]     io_axi_4_ar_bits_prot         ;
wire      [3:0]     io_axi_4_ar_bits_qos          ;
wire      [3:0]     io_axi_4_ar_bits_region       ;
wire      [2:0]     io_axi_4_ar_bits_size         ;
reg                 io_axi_4_w_ready              =0;
wire                io_axi_4_w_valid              ;
wire      [255:0]   io_axi_4_w_bits_data          ;
wire                io_axi_4_w_bits_last          ;
wire      [31:0]    io_axi_4_w_bits_strb          ;
wire                io_axi_4_r_ready              ;
reg                 io_axi_4_r_valid              =0;
reg       [255:0]   io_axi_4_r_bits_data          =0;
reg                 io_axi_4_r_bits_last          =0;
reg       [1:0]     io_axi_4_r_bits_resp          =0;
reg       [5:0]     io_axi_4_r_bits_id            =0;
wire                io_axi_4_b_ready              ;
reg                 io_axi_4_b_valid              =0;
reg       [5:0]     io_axi_4_b_bits_id            =0;
reg       [1:0]     io_axi_4_b_bits_resp          =0;
reg                 io_axi_5_aw_ready             =0;
wire                io_axi_5_aw_valid             ;
wire      [32:0]    io_axi_5_aw_bits_addr         ;
wire      [1:0]     io_axi_5_aw_bits_burst        ;
wire      [3:0]     io_axi_5_aw_bits_cache        ;
wire      [5:0]     io_axi_5_aw_bits_id           ;
wire      [3:0]     io_axi_5_aw_bits_len          ;
wire                io_axi_5_aw_bits_lock         ;
wire      [2:0]     io_axi_5_aw_bits_prot         ;
wire      [3:0]     io_axi_5_aw_bits_qos          ;
wire      [3:0]     io_axi_5_aw_bits_region       ;
wire      [2:0]     io_axi_5_aw_bits_size         ;
reg                 io_axi_5_ar_ready             =0;
wire                io_axi_5_ar_valid             ;
wire      [32:0]    io_axi_5_ar_bits_addr         ;
wire      [1:0]     io_axi_5_ar_bits_burst        ;
wire      [3:0]     io_axi_5_ar_bits_cache        ;
wire      [5:0]     io_axi_5_ar_bits_id           ;
wire      [3:0]     io_axi_5_ar_bits_len          ;
wire                io_axi_5_ar_bits_lock         ;
wire      [2:0]     io_axi_5_ar_bits_prot         ;
wire      [3:0]     io_axi_5_ar_bits_qos          ;
wire      [3:0]     io_axi_5_ar_bits_region       ;
wire      [2:0]     io_axi_5_ar_bits_size         ;
reg                 io_axi_5_w_ready              =0;
wire                io_axi_5_w_valid              ;
wire      [255:0]   io_axi_5_w_bits_data          ;
wire                io_axi_5_w_bits_last          ;
wire      [31:0]    io_axi_5_w_bits_strb          ;
wire                io_axi_5_r_ready              ;
reg                 io_axi_5_r_valid              =0;
reg       [255:0]   io_axi_5_r_bits_data          =0;
reg                 io_axi_5_r_bits_last          =0;
reg       [1:0]     io_axi_5_r_bits_resp          =0;
reg       [5:0]     io_axi_5_r_bits_id            =0;
wire                io_axi_5_b_ready              ;
reg                 io_axi_5_b_valid              =0;
reg       [5:0]     io_axi_5_b_bits_id            =0;
reg       [1:0]     io_axi_5_b_bits_resp          =0;
reg                 io_axi_6_aw_ready             =0;
wire                io_axi_6_aw_valid             ;
wire      [32:0]    io_axi_6_aw_bits_addr         ;
wire      [1:0]     io_axi_6_aw_bits_burst        ;
wire      [3:0]     io_axi_6_aw_bits_cache        ;
wire      [5:0]     io_axi_6_aw_bits_id           ;
wire      [3:0]     io_axi_6_aw_bits_len          ;
wire                io_axi_6_aw_bits_lock         ;
wire      [2:0]     io_axi_6_aw_bits_prot         ;
wire      [3:0]     io_axi_6_aw_bits_qos          ;
wire      [3:0]     io_axi_6_aw_bits_region       ;
wire      [2:0]     io_axi_6_aw_bits_size         ;
reg                 io_axi_6_ar_ready             =0;
wire                io_axi_6_ar_valid             ;
wire      [32:0]    io_axi_6_ar_bits_addr         ;
wire      [1:0]     io_axi_6_ar_bits_burst        ;
wire      [3:0]     io_axi_6_ar_bits_cache        ;
wire      [5:0]     io_axi_6_ar_bits_id           ;
wire      [3:0]     io_axi_6_ar_bits_len          ;
wire                io_axi_6_ar_bits_lock         ;
wire      [2:0]     io_axi_6_ar_bits_prot         ;
wire      [3:0]     io_axi_6_ar_bits_qos          ;
wire      [3:0]     io_axi_6_ar_bits_region       ;
wire      [2:0]     io_axi_6_ar_bits_size         ;
reg                 io_axi_6_w_ready              =0;
wire                io_axi_6_w_valid              ;
wire      [255:0]   io_axi_6_w_bits_data          ;
wire                io_axi_6_w_bits_last          ;
wire      [31:0]    io_axi_6_w_bits_strb          ;
wire                io_axi_6_r_ready              ;
reg                 io_axi_6_r_valid              =0;
reg       [255:0]   io_axi_6_r_bits_data          =0;
reg                 io_axi_6_r_bits_last          =0;
reg       [1:0]     io_axi_6_r_bits_resp          =0;
reg       [5:0]     io_axi_6_r_bits_id            =0;
wire                io_axi_6_b_ready              ;
reg                 io_axi_6_b_valid              =0;
reg       [5:0]     io_axi_6_b_bits_id            =0;
reg       [1:0]     io_axi_6_b_bits_resp          =0;
reg                 io_axi_7_aw_ready             =0;
wire                io_axi_7_aw_valid             ;
wire      [32:0]    io_axi_7_aw_bits_addr         ;
wire      [1:0]     io_axi_7_aw_bits_burst        ;
wire      [3:0]     io_axi_7_aw_bits_cache        ;
wire      [5:0]     io_axi_7_aw_bits_id           ;
wire      [3:0]     io_axi_7_aw_bits_len          ;
wire                io_axi_7_aw_bits_lock         ;
wire      [2:0]     io_axi_7_aw_bits_prot         ;
wire      [3:0]     io_axi_7_aw_bits_qos          ;
wire      [3:0]     io_axi_7_aw_bits_region       ;
wire      [2:0]     io_axi_7_aw_bits_size         ;
reg                 io_axi_7_ar_ready             =0;
wire                io_axi_7_ar_valid             ;
wire      [32:0]    io_axi_7_ar_bits_addr         ;
wire      [1:0]     io_axi_7_ar_bits_burst        ;
wire      [3:0]     io_axi_7_ar_bits_cache        ;
wire      [5:0]     io_axi_7_ar_bits_id           ;
wire      [3:0]     io_axi_7_ar_bits_len          ;
wire                io_axi_7_ar_bits_lock         ;
wire      [2:0]     io_axi_7_ar_bits_prot         ;
wire      [3:0]     io_axi_7_ar_bits_qos          ;
wire      [3:0]     io_axi_7_ar_bits_region       ;
wire      [2:0]     io_axi_7_ar_bits_size         ;
reg                 io_axi_7_w_ready              =0;
wire                io_axi_7_w_valid              ;
wire      [255:0]   io_axi_7_w_bits_data          ;
wire                io_axi_7_w_bits_last          ;
wire      [31:0]    io_axi_7_w_bits_strb          ;
wire                io_axi_7_r_ready              ;
reg                 io_axi_7_r_valid              =0;
reg       [255:0]   io_axi_7_r_bits_data          =0;
reg                 io_axi_7_r_bits_last          =0;
reg       [1:0]     io_axi_7_r_bits_resp          =0;
reg       [5:0]     io_axi_7_r_bits_id            =0;
wire                io_axi_7_b_ready              ;
reg                 io_axi_7_b_valid              =0;
reg       [5:0]     io_axi_7_b_bits_id            =0;
reg       [1:0]     io_axi_7_b_bits_resp          =0;
reg                 io_axi_8_aw_ready             =0;
wire                io_axi_8_aw_valid             ;
wire      [32:0]    io_axi_8_aw_bits_addr         ;
wire      [1:0]     io_axi_8_aw_bits_burst        ;
wire      [3:0]     io_axi_8_aw_bits_cache        ;
wire      [5:0]     io_axi_8_aw_bits_id           ;
wire      [3:0]     io_axi_8_aw_bits_len          ;
wire                io_axi_8_aw_bits_lock         ;
wire      [2:0]     io_axi_8_aw_bits_prot         ;
wire      [3:0]     io_axi_8_aw_bits_qos          ;
wire      [3:0]     io_axi_8_aw_bits_region       ;
wire      [2:0]     io_axi_8_aw_bits_size         ;
reg                 io_axi_8_ar_ready             =0;
wire                io_axi_8_ar_valid             ;
wire      [32:0]    io_axi_8_ar_bits_addr         ;
wire      [1:0]     io_axi_8_ar_bits_burst        ;
wire      [3:0]     io_axi_8_ar_bits_cache        ;
wire      [5:0]     io_axi_8_ar_bits_id           ;
wire      [3:0]     io_axi_8_ar_bits_len          ;
wire                io_axi_8_ar_bits_lock         ;
wire      [2:0]     io_axi_8_ar_bits_prot         ;
wire      [3:0]     io_axi_8_ar_bits_qos          ;
wire      [3:0]     io_axi_8_ar_bits_region       ;
wire      [2:0]     io_axi_8_ar_bits_size         ;
reg                 io_axi_8_w_ready              =0;
wire                io_axi_8_w_valid              ;
wire      [255:0]   io_axi_8_w_bits_data          ;
wire                io_axi_8_w_bits_last          ;
wire      [31:0]    io_axi_8_w_bits_strb          ;
wire                io_axi_8_r_ready              ;
reg                 io_axi_8_r_valid              =0;
reg       [255:0]   io_axi_8_r_bits_data          =0;
reg                 io_axi_8_r_bits_last          =0;
reg       [1:0]     io_axi_8_r_bits_resp          =0;
reg       [5:0]     io_axi_8_r_bits_id            =0;
wire                io_axi_8_b_ready              ;
reg                 io_axi_8_b_valid              =0;
reg       [5:0]     io_axi_8_b_bits_id            =0;
reg       [1:0]     io_axi_8_b_bits_resp          =0;
reg                 io_axi_9_aw_ready             =0;
wire                io_axi_9_aw_valid             ;
wire      [32:0]    io_axi_9_aw_bits_addr         ;
wire      [1:0]     io_axi_9_aw_bits_burst        ;
wire      [3:0]     io_axi_9_aw_bits_cache        ;
wire      [5:0]     io_axi_9_aw_bits_id           ;
wire      [3:0]     io_axi_9_aw_bits_len          ;
wire                io_axi_9_aw_bits_lock         ;
wire      [2:0]     io_axi_9_aw_bits_prot         ;
wire      [3:0]     io_axi_9_aw_bits_qos          ;
wire      [3:0]     io_axi_9_aw_bits_region       ;
wire      [2:0]     io_axi_9_aw_bits_size         ;
reg                 io_axi_9_ar_ready             =0;
wire                io_axi_9_ar_valid             ;
wire      [32:0]    io_axi_9_ar_bits_addr         ;
wire      [1:0]     io_axi_9_ar_bits_burst        ;
wire      [3:0]     io_axi_9_ar_bits_cache        ;
wire      [5:0]     io_axi_9_ar_bits_id           ;
wire      [3:0]     io_axi_9_ar_bits_len          ;
wire                io_axi_9_ar_bits_lock         ;
wire      [2:0]     io_axi_9_ar_bits_prot         ;
wire      [3:0]     io_axi_9_ar_bits_qos          ;
wire      [3:0]     io_axi_9_ar_bits_region       ;
wire      [2:0]     io_axi_9_ar_bits_size         ;
reg                 io_axi_9_w_ready              =0;
wire                io_axi_9_w_valid              ;
wire      [255:0]   io_axi_9_w_bits_data          ;
wire                io_axi_9_w_bits_last          ;
wire      [31:0]    io_axi_9_w_bits_strb          ;
wire                io_axi_9_r_ready              ;
reg                 io_axi_9_r_valid              =0;
reg       [255:0]   io_axi_9_r_bits_data          =0;
reg                 io_axi_9_r_bits_last          =0;
reg       [1:0]     io_axi_9_r_bits_resp          =0;
reg       [5:0]     io_axi_9_r_bits_id            =0;
wire                io_axi_9_b_ready              ;
reg                 io_axi_9_b_valid              =0;
reg       [5:0]     io_axi_9_b_bits_id            =0;
reg       [1:0]     io_axi_9_b_bits_resp          =0;
reg                 io_axi_10_aw_ready            =0;
wire                io_axi_10_aw_valid            ;
wire      [32:0]    io_axi_10_aw_bits_addr        ;
wire      [1:0]     io_axi_10_aw_bits_burst       ;
wire      [3:0]     io_axi_10_aw_bits_cache       ;
wire      [5:0]     io_axi_10_aw_bits_id          ;
wire      [3:0]     io_axi_10_aw_bits_len         ;
wire                io_axi_10_aw_bits_lock        ;
wire      [2:0]     io_axi_10_aw_bits_prot        ;
wire      [3:0]     io_axi_10_aw_bits_qos         ;
wire      [3:0]     io_axi_10_aw_bits_region      ;
wire      [2:0]     io_axi_10_aw_bits_size        ;
reg                 io_axi_10_ar_ready            =0;
wire                io_axi_10_ar_valid            ;
wire      [32:0]    io_axi_10_ar_bits_addr        ;
wire      [1:0]     io_axi_10_ar_bits_burst       ;
wire      [3:0]     io_axi_10_ar_bits_cache       ;
wire      [5:0]     io_axi_10_ar_bits_id          ;
wire      [3:0]     io_axi_10_ar_bits_len         ;
wire                io_axi_10_ar_bits_lock        ;
wire      [2:0]     io_axi_10_ar_bits_prot        ;
wire      [3:0]     io_axi_10_ar_bits_qos         ;
wire      [3:0]     io_axi_10_ar_bits_region      ;
wire      [2:0]     io_axi_10_ar_bits_size        ;
reg                 io_axi_10_w_ready             =0;
wire                io_axi_10_w_valid             ;
wire      [255:0]   io_axi_10_w_bits_data         ;
wire                io_axi_10_w_bits_last         ;
wire      [31:0]    io_axi_10_w_bits_strb         ;
wire                io_axi_10_r_ready             ;
reg                 io_axi_10_r_valid             =0;
reg       [255:0]   io_axi_10_r_bits_data         =0;
reg                 io_axi_10_r_bits_last         =0;
reg       [1:0]     io_axi_10_r_bits_resp         =0;
reg       [5:0]     io_axi_10_r_bits_id           =0;
wire                io_axi_10_b_ready             ;
reg                 io_axi_10_b_valid             =0;
reg       [5:0]     io_axi_10_b_bits_id           =0;
reg       [1:0]     io_axi_10_b_bits_resp         =0;
reg                 io_axi_11_aw_ready            =0;
wire                io_axi_11_aw_valid            ;
wire      [32:0]    io_axi_11_aw_bits_addr        ;
wire      [1:0]     io_axi_11_aw_bits_burst       ;
wire      [3:0]     io_axi_11_aw_bits_cache       ;
wire      [5:0]     io_axi_11_aw_bits_id          ;
wire      [3:0]     io_axi_11_aw_bits_len         ;
wire                io_axi_11_aw_bits_lock        ;
wire      [2:0]     io_axi_11_aw_bits_prot        ;
wire      [3:0]     io_axi_11_aw_bits_qos         ;
wire      [3:0]     io_axi_11_aw_bits_region      ;
wire      [2:0]     io_axi_11_aw_bits_size        ;
reg                 io_axi_11_ar_ready            =0;
wire                io_axi_11_ar_valid            ;
wire      [32:0]    io_axi_11_ar_bits_addr        ;
wire      [1:0]     io_axi_11_ar_bits_burst       ;
wire      [3:0]     io_axi_11_ar_bits_cache       ;
wire      [5:0]     io_axi_11_ar_bits_id          ;
wire      [3:0]     io_axi_11_ar_bits_len         ;
wire                io_axi_11_ar_bits_lock        ;
wire      [2:0]     io_axi_11_ar_bits_prot        ;
wire      [3:0]     io_axi_11_ar_bits_qos         ;
wire      [3:0]     io_axi_11_ar_bits_region      ;
wire      [2:0]     io_axi_11_ar_bits_size        ;
reg                 io_axi_11_w_ready             =0;
wire                io_axi_11_w_valid             ;
wire      [255:0]   io_axi_11_w_bits_data         ;
wire                io_axi_11_w_bits_last         ;
wire      [31:0]    io_axi_11_w_bits_strb         ;
wire                io_axi_11_r_ready             ;
reg                 io_axi_11_r_valid             =0;
reg       [255:0]   io_axi_11_r_bits_data         =0;
reg                 io_axi_11_r_bits_last         =0;
reg       [1:0]     io_axi_11_r_bits_resp         =0;
reg       [5:0]     io_axi_11_r_bits_id           =0;
wire                io_axi_11_b_ready             ;
reg                 io_axi_11_b_valid             =0;
reg       [5:0]     io_axi_11_b_bits_id           =0;
reg       [1:0]     io_axi_11_b_bits_resp         =0;
reg                 io_axi_12_aw_ready            =0;
wire                io_axi_12_aw_valid            ;
wire      [32:0]    io_axi_12_aw_bits_addr        ;
wire      [1:0]     io_axi_12_aw_bits_burst       ;
wire      [3:0]     io_axi_12_aw_bits_cache       ;
wire      [5:0]     io_axi_12_aw_bits_id          ;
wire      [3:0]     io_axi_12_aw_bits_len         ;
wire                io_axi_12_aw_bits_lock        ;
wire      [2:0]     io_axi_12_aw_bits_prot        ;
wire      [3:0]     io_axi_12_aw_bits_qos         ;
wire      [3:0]     io_axi_12_aw_bits_region      ;
wire      [2:0]     io_axi_12_aw_bits_size        ;
reg                 io_axi_12_ar_ready            =0;
wire                io_axi_12_ar_valid            ;
wire      [32:0]    io_axi_12_ar_bits_addr        ;
wire      [1:0]     io_axi_12_ar_bits_burst       ;
wire      [3:0]     io_axi_12_ar_bits_cache       ;
wire      [5:0]     io_axi_12_ar_bits_id          ;
wire      [3:0]     io_axi_12_ar_bits_len         ;
wire                io_axi_12_ar_bits_lock        ;
wire      [2:0]     io_axi_12_ar_bits_prot        ;
wire      [3:0]     io_axi_12_ar_bits_qos         ;
wire      [3:0]     io_axi_12_ar_bits_region      ;
wire      [2:0]     io_axi_12_ar_bits_size        ;
reg                 io_axi_12_w_ready             =0;
wire                io_axi_12_w_valid             ;
wire      [255:0]   io_axi_12_w_bits_data         ;
wire                io_axi_12_w_bits_last         ;
wire      [31:0]    io_axi_12_w_bits_strb         ;
wire                io_axi_12_r_ready             ;
reg                 io_axi_12_r_valid             =0;
reg       [255:0]   io_axi_12_r_bits_data         =0;
reg                 io_axi_12_r_bits_last         =0;
reg       [1:0]     io_axi_12_r_bits_resp         =0;
reg       [5:0]     io_axi_12_r_bits_id           =0;
wire                io_axi_12_b_ready             ;
reg                 io_axi_12_b_valid             =0;
reg       [5:0]     io_axi_12_b_bits_id           =0;
reg       [1:0]     io_axi_12_b_bits_resp         =0;
reg                 io_axi_13_aw_ready            =0;
wire                io_axi_13_aw_valid            ;
wire      [32:0]    io_axi_13_aw_bits_addr        ;
wire      [1:0]     io_axi_13_aw_bits_burst       ;
wire      [3:0]     io_axi_13_aw_bits_cache       ;
wire      [5:0]     io_axi_13_aw_bits_id          ;
wire      [3:0]     io_axi_13_aw_bits_len         ;
wire                io_axi_13_aw_bits_lock        ;
wire      [2:0]     io_axi_13_aw_bits_prot        ;
wire      [3:0]     io_axi_13_aw_bits_qos         ;
wire      [3:0]     io_axi_13_aw_bits_region      ;
wire      [2:0]     io_axi_13_aw_bits_size        ;
reg                 io_axi_13_ar_ready            =0;
wire                io_axi_13_ar_valid            ;
wire      [32:0]    io_axi_13_ar_bits_addr        ;
wire      [1:0]     io_axi_13_ar_bits_burst       ;
wire      [3:0]     io_axi_13_ar_bits_cache       ;
wire      [5:0]     io_axi_13_ar_bits_id          ;
wire      [3:0]     io_axi_13_ar_bits_len         ;
wire                io_axi_13_ar_bits_lock        ;
wire      [2:0]     io_axi_13_ar_bits_prot        ;
wire      [3:0]     io_axi_13_ar_bits_qos         ;
wire      [3:0]     io_axi_13_ar_bits_region      ;
wire      [2:0]     io_axi_13_ar_bits_size        ;
reg                 io_axi_13_w_ready             =0;
wire                io_axi_13_w_valid             ;
wire      [255:0]   io_axi_13_w_bits_data         ;
wire                io_axi_13_w_bits_last         ;
wire      [31:0]    io_axi_13_w_bits_strb         ;
wire                io_axi_13_r_ready             ;
reg                 io_axi_13_r_valid             =0;
reg       [255:0]   io_axi_13_r_bits_data         =0;
reg                 io_axi_13_r_bits_last         =0;
reg       [1:0]     io_axi_13_r_bits_resp         =0;
reg       [5:0]     io_axi_13_r_bits_id           =0;
wire                io_axi_13_b_ready             ;
reg                 io_axi_13_b_valid             =0;
reg       [5:0]     io_axi_13_b_bits_id           =0;
reg       [1:0]     io_axi_13_b_bits_resp         =0;
reg                 io_axi_14_aw_ready            =0;
wire                io_axi_14_aw_valid            ;
wire      [32:0]    io_axi_14_aw_bits_addr        ;
wire      [1:0]     io_axi_14_aw_bits_burst       ;
wire      [3:0]     io_axi_14_aw_bits_cache       ;
wire      [5:0]     io_axi_14_aw_bits_id          ;
wire      [3:0]     io_axi_14_aw_bits_len         ;
wire                io_axi_14_aw_bits_lock        ;
wire      [2:0]     io_axi_14_aw_bits_prot        ;
wire      [3:0]     io_axi_14_aw_bits_qos         ;
wire      [3:0]     io_axi_14_aw_bits_region      ;
wire      [2:0]     io_axi_14_aw_bits_size        ;
reg                 io_axi_14_ar_ready            =0;
wire                io_axi_14_ar_valid            ;
wire      [32:0]    io_axi_14_ar_bits_addr        ;
wire      [1:0]     io_axi_14_ar_bits_burst       ;
wire      [3:0]     io_axi_14_ar_bits_cache       ;
wire      [5:0]     io_axi_14_ar_bits_id          ;
wire      [3:0]     io_axi_14_ar_bits_len         ;
wire                io_axi_14_ar_bits_lock        ;
wire      [2:0]     io_axi_14_ar_bits_prot        ;
wire      [3:0]     io_axi_14_ar_bits_qos         ;
wire      [3:0]     io_axi_14_ar_bits_region      ;
wire      [2:0]     io_axi_14_ar_bits_size        ;
reg                 io_axi_14_w_ready             =0;
wire                io_axi_14_w_valid             ;
wire      [255:0]   io_axi_14_w_bits_data         ;
wire                io_axi_14_w_bits_last         ;
wire      [31:0]    io_axi_14_w_bits_strb         ;
wire                io_axi_14_r_ready             ;
reg                 io_axi_14_r_valid             =0;
reg       [255:0]   io_axi_14_r_bits_data         =0;
reg                 io_axi_14_r_bits_last         =0;
reg       [1:0]     io_axi_14_r_bits_resp         =0;
reg       [5:0]     io_axi_14_r_bits_id           =0;
wire                io_axi_14_b_ready             ;
reg                 io_axi_14_b_valid             =0;
reg       [5:0]     io_axi_14_b_bits_id           =0;
reg       [1:0]     io_axi_14_b_bits_resp         =0;
reg                 io_axi_15_aw_ready            =0;
wire                io_axi_15_aw_valid            ;
wire      [32:0]    io_axi_15_aw_bits_addr        ;
wire      [1:0]     io_axi_15_aw_bits_burst       ;
wire      [3:0]     io_axi_15_aw_bits_cache       ;
wire      [5:0]     io_axi_15_aw_bits_id          ;
wire      [3:0]     io_axi_15_aw_bits_len         ;
wire                io_axi_15_aw_bits_lock        ;
wire      [2:0]     io_axi_15_aw_bits_prot        ;
wire      [3:0]     io_axi_15_aw_bits_qos         ;
wire      [3:0]     io_axi_15_aw_bits_region      ;
wire      [2:0]     io_axi_15_aw_bits_size        ;
reg                 io_axi_15_ar_ready            =0;
wire                io_axi_15_ar_valid            ;
wire      [32:0]    io_axi_15_ar_bits_addr        ;
wire      [1:0]     io_axi_15_ar_bits_burst       ;
wire      [3:0]     io_axi_15_ar_bits_cache       ;
wire      [5:0]     io_axi_15_ar_bits_id          ;
wire      [3:0]     io_axi_15_ar_bits_len         ;
wire                io_axi_15_ar_bits_lock        ;
wire      [2:0]     io_axi_15_ar_bits_prot        ;
wire      [3:0]     io_axi_15_ar_bits_qos         ;
wire      [3:0]     io_axi_15_ar_bits_region      ;
wire      [2:0]     io_axi_15_ar_bits_size        ;
reg                 io_axi_15_w_ready             =0;
wire                io_axi_15_w_valid             ;
wire      [255:0]   io_axi_15_w_bits_data         ;
wire                io_axi_15_w_bits_last         ;
wire      [31:0]    io_axi_15_w_bits_strb         ;
wire                io_axi_15_r_ready             ;
reg                 io_axi_15_r_valid             =0;
reg       [255:0]   io_axi_15_r_bits_data         =0;
reg                 io_axi_15_r_bits_last         =0;
reg       [1:0]     io_axi_15_r_bits_resp         =0;
reg       [5:0]     io_axi_15_r_bits_id           =0;
wire                io_axi_15_b_ready             ;
reg                 io_axi_15_b_valid             =0;
reg       [5:0]     io_axi_15_b_bits_id           =0;
reg       [1:0]     io_axi_15_b_bits_resp         =0;
reg                 io_axi_16_aw_ready            =0;
wire                io_axi_16_aw_valid            ;
wire      [32:0]    io_axi_16_aw_bits_addr        ;
wire      [1:0]     io_axi_16_aw_bits_burst       ;
wire      [3:0]     io_axi_16_aw_bits_cache       ;
wire      [5:0]     io_axi_16_aw_bits_id          ;
wire      [3:0]     io_axi_16_aw_bits_len         ;
wire                io_axi_16_aw_bits_lock        ;
wire      [2:0]     io_axi_16_aw_bits_prot        ;
wire      [3:0]     io_axi_16_aw_bits_qos         ;
wire      [3:0]     io_axi_16_aw_bits_region      ;
wire      [2:0]     io_axi_16_aw_bits_size        ;
reg                 io_axi_16_ar_ready            =0;
wire                io_axi_16_ar_valid            ;
wire      [32:0]    io_axi_16_ar_bits_addr        ;
wire      [1:0]     io_axi_16_ar_bits_burst       ;
wire      [3:0]     io_axi_16_ar_bits_cache       ;
wire      [5:0]     io_axi_16_ar_bits_id          ;
wire      [3:0]     io_axi_16_ar_bits_len         ;
wire                io_axi_16_ar_bits_lock        ;
wire      [2:0]     io_axi_16_ar_bits_prot        ;
wire      [3:0]     io_axi_16_ar_bits_qos         ;
wire      [3:0]     io_axi_16_ar_bits_region      ;
wire      [2:0]     io_axi_16_ar_bits_size        ;
reg                 io_axi_16_w_ready             =0;
wire                io_axi_16_w_valid             ;
wire      [255:0]   io_axi_16_w_bits_data         ;
wire                io_axi_16_w_bits_last         ;
wire      [31:0]    io_axi_16_w_bits_strb         ;
wire                io_axi_16_r_ready             ;
reg                 io_axi_16_r_valid             =0;
reg       [255:0]   io_axi_16_r_bits_data         =0;
reg                 io_axi_16_r_bits_last         =0;
reg       [1:0]     io_axi_16_r_bits_resp         =0;
reg       [5:0]     io_axi_16_r_bits_id           =0;
wire                io_axi_16_b_ready             ;
reg                 io_axi_16_b_valid             =0;
reg       [5:0]     io_axi_16_b_bits_id           =0;
reg       [1:0]     io_axi_16_b_bits_resp         =0;
reg                 io_axi_17_aw_ready            =0;
wire                io_axi_17_aw_valid            ;
wire      [32:0]    io_axi_17_aw_bits_addr        ;
wire      [1:0]     io_axi_17_aw_bits_burst       ;
wire      [3:0]     io_axi_17_aw_bits_cache       ;
wire      [5:0]     io_axi_17_aw_bits_id          ;
wire      [3:0]     io_axi_17_aw_bits_len         ;
wire                io_axi_17_aw_bits_lock        ;
wire      [2:0]     io_axi_17_aw_bits_prot        ;
wire      [3:0]     io_axi_17_aw_bits_qos         ;
wire      [3:0]     io_axi_17_aw_bits_region      ;
wire      [2:0]     io_axi_17_aw_bits_size        ;
reg                 io_axi_17_ar_ready            =0;
wire                io_axi_17_ar_valid            ;
wire      [32:0]    io_axi_17_ar_bits_addr        ;
wire      [1:0]     io_axi_17_ar_bits_burst       ;
wire      [3:0]     io_axi_17_ar_bits_cache       ;
wire      [5:0]     io_axi_17_ar_bits_id          ;
wire      [3:0]     io_axi_17_ar_bits_len         ;
wire                io_axi_17_ar_bits_lock        ;
wire      [2:0]     io_axi_17_ar_bits_prot        ;
wire      [3:0]     io_axi_17_ar_bits_qos         ;
wire      [3:0]     io_axi_17_ar_bits_region      ;
wire      [2:0]     io_axi_17_ar_bits_size        ;
reg                 io_axi_17_w_ready             =0;
wire                io_axi_17_w_valid             ;
wire      [255:0]   io_axi_17_w_bits_data         ;
wire                io_axi_17_w_bits_last         ;
wire      [31:0]    io_axi_17_w_bits_strb         ;
wire                io_axi_17_r_ready             ;
reg                 io_axi_17_r_valid             =0;
reg       [255:0]   io_axi_17_r_bits_data         =0;
reg                 io_axi_17_r_bits_last         =0;
reg       [1:0]     io_axi_17_r_bits_resp         =0;
reg       [5:0]     io_axi_17_r_bits_id           =0;
wire                io_axi_17_b_ready             ;
reg                 io_axi_17_b_valid             =0;
reg       [5:0]     io_axi_17_b_bits_id           =0;
reg       [1:0]     io_axi_17_b_bits_resp         =0;
reg                 io_axi_18_aw_ready            =0;
wire                io_axi_18_aw_valid            ;
wire      [32:0]    io_axi_18_aw_bits_addr        ;
wire      [1:0]     io_axi_18_aw_bits_burst       ;
wire      [3:0]     io_axi_18_aw_bits_cache       ;
wire      [5:0]     io_axi_18_aw_bits_id          ;
wire      [3:0]     io_axi_18_aw_bits_len         ;
wire                io_axi_18_aw_bits_lock        ;
wire      [2:0]     io_axi_18_aw_bits_prot        ;
wire      [3:0]     io_axi_18_aw_bits_qos         ;
wire      [3:0]     io_axi_18_aw_bits_region      ;
wire      [2:0]     io_axi_18_aw_bits_size        ;
reg                 io_axi_18_ar_ready            =0;
wire                io_axi_18_ar_valid            ;
wire      [32:0]    io_axi_18_ar_bits_addr        ;
wire      [1:0]     io_axi_18_ar_bits_burst       ;
wire      [3:0]     io_axi_18_ar_bits_cache       ;
wire      [5:0]     io_axi_18_ar_bits_id          ;
wire      [3:0]     io_axi_18_ar_bits_len         ;
wire                io_axi_18_ar_bits_lock        ;
wire      [2:0]     io_axi_18_ar_bits_prot        ;
wire      [3:0]     io_axi_18_ar_bits_qos         ;
wire      [3:0]     io_axi_18_ar_bits_region      ;
wire      [2:0]     io_axi_18_ar_bits_size        ;
reg                 io_axi_18_w_ready             =0;
wire                io_axi_18_w_valid             ;
wire      [255:0]   io_axi_18_w_bits_data         ;
wire                io_axi_18_w_bits_last         ;
wire      [31:0]    io_axi_18_w_bits_strb         ;
wire                io_axi_18_r_ready             ;
reg                 io_axi_18_r_valid             =0;
reg       [255:0]   io_axi_18_r_bits_data         =0;
reg                 io_axi_18_r_bits_last         =0;
reg       [1:0]     io_axi_18_r_bits_resp         =0;
reg       [5:0]     io_axi_18_r_bits_id           =0;
wire                io_axi_18_b_ready             ;
reg                 io_axi_18_b_valid             =0;
reg       [5:0]     io_axi_18_b_bits_id           =0;
reg       [1:0]     io_axi_18_b_bits_resp         =0;
reg                 io_axi_19_aw_ready            =0;
wire                io_axi_19_aw_valid            ;
wire      [32:0]    io_axi_19_aw_bits_addr        ;
wire      [1:0]     io_axi_19_aw_bits_burst       ;
wire      [3:0]     io_axi_19_aw_bits_cache       ;
wire      [5:0]     io_axi_19_aw_bits_id          ;
wire      [3:0]     io_axi_19_aw_bits_len         ;
wire                io_axi_19_aw_bits_lock        ;
wire      [2:0]     io_axi_19_aw_bits_prot        ;
wire      [3:0]     io_axi_19_aw_bits_qos         ;
wire      [3:0]     io_axi_19_aw_bits_region      ;
wire      [2:0]     io_axi_19_aw_bits_size        ;
reg                 io_axi_19_ar_ready            =0;
wire                io_axi_19_ar_valid            ;
wire      [32:0]    io_axi_19_ar_bits_addr        ;
wire      [1:0]     io_axi_19_ar_bits_burst       ;
wire      [3:0]     io_axi_19_ar_bits_cache       ;
wire      [5:0]     io_axi_19_ar_bits_id          ;
wire      [3:0]     io_axi_19_ar_bits_len         ;
wire                io_axi_19_ar_bits_lock        ;
wire      [2:0]     io_axi_19_ar_bits_prot        ;
wire      [3:0]     io_axi_19_ar_bits_qos         ;
wire      [3:0]     io_axi_19_ar_bits_region      ;
wire      [2:0]     io_axi_19_ar_bits_size        ;
reg                 io_axi_19_w_ready             =0;
wire                io_axi_19_w_valid             ;
wire      [255:0]   io_axi_19_w_bits_data         ;
wire                io_axi_19_w_bits_last         ;
wire      [31:0]    io_axi_19_w_bits_strb         ;
wire                io_axi_19_r_ready             ;
reg                 io_axi_19_r_valid             =0;
reg       [255:0]   io_axi_19_r_bits_data         =0;
reg                 io_axi_19_r_bits_last         =0;
reg       [1:0]     io_axi_19_r_bits_resp         =0;
reg       [5:0]     io_axi_19_r_bits_id           =0;
wire                io_axi_19_b_ready             ;
reg                 io_axi_19_b_valid             =0;
reg       [5:0]     io_axi_19_b_bits_id           =0;
reg       [1:0]     io_axi_19_b_bits_resp         =0;
reg                 io_axi_20_aw_ready            =0;
wire                io_axi_20_aw_valid            ;
wire      [32:0]    io_axi_20_aw_bits_addr        ;
wire      [1:0]     io_axi_20_aw_bits_burst       ;
wire      [3:0]     io_axi_20_aw_bits_cache       ;
wire      [5:0]     io_axi_20_aw_bits_id          ;
wire      [3:0]     io_axi_20_aw_bits_len         ;
wire                io_axi_20_aw_bits_lock        ;
wire      [2:0]     io_axi_20_aw_bits_prot        ;
wire      [3:0]     io_axi_20_aw_bits_qos         ;
wire      [3:0]     io_axi_20_aw_bits_region      ;
wire      [2:0]     io_axi_20_aw_bits_size        ;
reg                 io_axi_20_ar_ready            =0;
wire                io_axi_20_ar_valid            ;
wire      [32:0]    io_axi_20_ar_bits_addr        ;
wire      [1:0]     io_axi_20_ar_bits_burst       ;
wire      [3:0]     io_axi_20_ar_bits_cache       ;
wire      [5:0]     io_axi_20_ar_bits_id          ;
wire      [3:0]     io_axi_20_ar_bits_len         ;
wire                io_axi_20_ar_bits_lock        ;
wire      [2:0]     io_axi_20_ar_bits_prot        ;
wire      [3:0]     io_axi_20_ar_bits_qos         ;
wire      [3:0]     io_axi_20_ar_bits_region      ;
wire      [2:0]     io_axi_20_ar_bits_size        ;
reg                 io_axi_20_w_ready             =0;
wire                io_axi_20_w_valid             ;
wire      [255:0]   io_axi_20_w_bits_data         ;
wire                io_axi_20_w_bits_last         ;
wire      [31:0]    io_axi_20_w_bits_strb         ;
wire                io_axi_20_r_ready             ;
reg                 io_axi_20_r_valid             =0;
reg       [255:0]   io_axi_20_r_bits_data         =0;
reg                 io_axi_20_r_bits_last         =0;
reg       [1:0]     io_axi_20_r_bits_resp         =0;
reg       [5:0]     io_axi_20_r_bits_id           =0;
wire                io_axi_20_b_ready             ;
reg                 io_axi_20_b_valid             =0;
reg       [5:0]     io_axi_20_b_bits_id           =0;
reg       [1:0]     io_axi_20_b_bits_resp         =0;
reg                 io_axi_21_aw_ready            =0;
wire                io_axi_21_aw_valid            ;
wire      [32:0]    io_axi_21_aw_bits_addr        ;
wire      [1:0]     io_axi_21_aw_bits_burst       ;
wire      [3:0]     io_axi_21_aw_bits_cache       ;
wire      [5:0]     io_axi_21_aw_bits_id          ;
wire      [3:0]     io_axi_21_aw_bits_len         ;
wire                io_axi_21_aw_bits_lock        ;
wire      [2:0]     io_axi_21_aw_bits_prot        ;
wire      [3:0]     io_axi_21_aw_bits_qos         ;
wire      [3:0]     io_axi_21_aw_bits_region      ;
wire      [2:0]     io_axi_21_aw_bits_size        ;
reg                 io_axi_21_ar_ready            =0;
wire                io_axi_21_ar_valid            ;
wire      [32:0]    io_axi_21_ar_bits_addr        ;
wire      [1:0]     io_axi_21_ar_bits_burst       ;
wire      [3:0]     io_axi_21_ar_bits_cache       ;
wire      [5:0]     io_axi_21_ar_bits_id          ;
wire      [3:0]     io_axi_21_ar_bits_len         ;
wire                io_axi_21_ar_bits_lock        ;
wire      [2:0]     io_axi_21_ar_bits_prot        ;
wire      [3:0]     io_axi_21_ar_bits_qos         ;
wire      [3:0]     io_axi_21_ar_bits_region      ;
wire      [2:0]     io_axi_21_ar_bits_size        ;
reg                 io_axi_21_w_ready             =0;
wire                io_axi_21_w_valid             ;
wire      [255:0]   io_axi_21_w_bits_data         ;
wire                io_axi_21_w_bits_last         ;
wire      [31:0]    io_axi_21_w_bits_strb         ;
wire                io_axi_21_r_ready             ;
reg                 io_axi_21_r_valid             =0;
reg       [255:0]   io_axi_21_r_bits_data         =0;
reg                 io_axi_21_r_bits_last         =0;
reg       [1:0]     io_axi_21_r_bits_resp         =0;
reg       [5:0]     io_axi_21_r_bits_id           =0;
wire                io_axi_21_b_ready             ;
reg                 io_axi_21_b_valid             =0;
reg       [5:0]     io_axi_21_b_bits_id           =0;
reg       [1:0]     io_axi_21_b_bits_resp         =0;
reg                 io_axi_22_aw_ready            =0;
wire                io_axi_22_aw_valid            ;
wire      [32:0]    io_axi_22_aw_bits_addr        ;
wire      [1:0]     io_axi_22_aw_bits_burst       ;
wire      [3:0]     io_axi_22_aw_bits_cache       ;
wire      [5:0]     io_axi_22_aw_bits_id          ;
wire      [3:0]     io_axi_22_aw_bits_len         ;
wire                io_axi_22_aw_bits_lock        ;
wire      [2:0]     io_axi_22_aw_bits_prot        ;
wire      [3:0]     io_axi_22_aw_bits_qos         ;
wire      [3:0]     io_axi_22_aw_bits_region      ;
wire      [2:0]     io_axi_22_aw_bits_size        ;
reg                 io_axi_22_ar_ready            =0;
wire                io_axi_22_ar_valid            ;
wire      [32:0]    io_axi_22_ar_bits_addr        ;
wire      [1:0]     io_axi_22_ar_bits_burst       ;
wire      [3:0]     io_axi_22_ar_bits_cache       ;
wire      [5:0]     io_axi_22_ar_bits_id          ;
wire      [3:0]     io_axi_22_ar_bits_len         ;
wire                io_axi_22_ar_bits_lock        ;
wire      [2:0]     io_axi_22_ar_bits_prot        ;
wire      [3:0]     io_axi_22_ar_bits_qos         ;
wire      [3:0]     io_axi_22_ar_bits_region      ;
wire      [2:0]     io_axi_22_ar_bits_size        ;
reg                 io_axi_22_w_ready             =0;
wire                io_axi_22_w_valid             ;
wire      [255:0]   io_axi_22_w_bits_data         ;
wire                io_axi_22_w_bits_last         ;
wire      [31:0]    io_axi_22_w_bits_strb         ;
wire                io_axi_22_r_ready             ;
reg                 io_axi_22_r_valid             =0;
reg       [255:0]   io_axi_22_r_bits_data         =0;
reg                 io_axi_22_r_bits_last         =0;
reg       [1:0]     io_axi_22_r_bits_resp         =0;
reg       [5:0]     io_axi_22_r_bits_id           =0;
wire                io_axi_22_b_ready             ;
reg                 io_axi_22_b_valid             =0;
reg       [5:0]     io_axi_22_b_bits_id           =0;
reg       [1:0]     io_axi_22_b_bits_resp         =0;
reg                 io_axi_23_aw_ready            =0;
wire                io_axi_23_aw_valid            ;
wire      [32:0]    io_axi_23_aw_bits_addr        ;
wire      [1:0]     io_axi_23_aw_bits_burst       ;
wire      [3:0]     io_axi_23_aw_bits_cache       ;
wire      [5:0]     io_axi_23_aw_bits_id          ;
wire      [3:0]     io_axi_23_aw_bits_len         ;
wire                io_axi_23_aw_bits_lock        ;
wire      [2:0]     io_axi_23_aw_bits_prot        ;
wire      [3:0]     io_axi_23_aw_bits_qos         ;
wire      [3:0]     io_axi_23_aw_bits_region      ;
wire      [2:0]     io_axi_23_aw_bits_size        ;
reg                 io_axi_23_ar_ready            =0;
wire                io_axi_23_ar_valid            ;
wire      [32:0]    io_axi_23_ar_bits_addr        ;
wire      [1:0]     io_axi_23_ar_bits_burst       ;
wire      [3:0]     io_axi_23_ar_bits_cache       ;
wire      [5:0]     io_axi_23_ar_bits_id          ;
wire      [3:0]     io_axi_23_ar_bits_len         ;
wire                io_axi_23_ar_bits_lock        ;
wire      [2:0]     io_axi_23_ar_bits_prot        ;
wire      [3:0]     io_axi_23_ar_bits_qos         ;
wire      [3:0]     io_axi_23_ar_bits_region      ;
wire      [2:0]     io_axi_23_ar_bits_size        ;
reg                 io_axi_23_w_ready             =0;
wire                io_axi_23_w_valid             ;
wire      [255:0]   io_axi_23_w_bits_data         ;
wire                io_axi_23_w_bits_last         ;
wire      [31:0]    io_axi_23_w_bits_strb         ;
wire                io_axi_23_r_ready             ;
reg                 io_axi_23_r_valid             =0;
reg       [255:0]   io_axi_23_r_bits_data         =0;
reg                 io_axi_23_r_bits_last         =0;
reg       [1:0]     io_axi_23_r_bits_resp         =0;
reg       [5:0]     io_axi_23_r_bits_id           =0;
wire                io_axi_23_b_ready             ;
reg                 io_axi_23_b_valid             =0;
reg       [5:0]     io_axi_23_b_bits_id           =0;
reg       [1:0]     io_axi_23_b_bits_resp         =0;
reg                 io_axi_24_aw_ready            =0;
wire                io_axi_24_aw_valid            ;
wire      [32:0]    io_axi_24_aw_bits_addr        ;
wire      [1:0]     io_axi_24_aw_bits_burst       ;
wire      [3:0]     io_axi_24_aw_bits_cache       ;
wire      [5:0]     io_axi_24_aw_bits_id          ;
wire      [3:0]     io_axi_24_aw_bits_len         ;
wire                io_axi_24_aw_bits_lock        ;
wire      [2:0]     io_axi_24_aw_bits_prot        ;
wire      [3:0]     io_axi_24_aw_bits_qos         ;
wire      [3:0]     io_axi_24_aw_bits_region      ;
wire      [2:0]     io_axi_24_aw_bits_size        ;
reg                 io_axi_24_ar_ready            =0;
wire                io_axi_24_ar_valid            ;
wire      [32:0]    io_axi_24_ar_bits_addr        ;
wire      [1:0]     io_axi_24_ar_bits_burst       ;
wire      [3:0]     io_axi_24_ar_bits_cache       ;
wire      [5:0]     io_axi_24_ar_bits_id          ;
wire      [3:0]     io_axi_24_ar_bits_len         ;
wire                io_axi_24_ar_bits_lock        ;
wire      [2:0]     io_axi_24_ar_bits_prot        ;
wire      [3:0]     io_axi_24_ar_bits_qos         ;
wire      [3:0]     io_axi_24_ar_bits_region      ;
wire      [2:0]     io_axi_24_ar_bits_size        ;
reg                 io_axi_24_w_ready             =0;
wire                io_axi_24_w_valid             ;
wire      [255:0]   io_axi_24_w_bits_data         ;
wire                io_axi_24_w_bits_last         ;
wire      [31:0]    io_axi_24_w_bits_strb         ;
wire                io_axi_24_r_ready             ;
reg                 io_axi_24_r_valid             =0;
reg       [255:0]   io_axi_24_r_bits_data         =0;
reg                 io_axi_24_r_bits_last         =0;
reg       [1:0]     io_axi_24_r_bits_resp         =0;
reg       [5:0]     io_axi_24_r_bits_id           =0;
wire                io_axi_24_b_ready             ;
reg                 io_axi_24_b_valid             =0;
reg       [5:0]     io_axi_24_b_bits_id           =0;
reg       [1:0]     io_axi_24_b_bits_resp         =0;
reg                 io_axi_25_aw_ready            =0;
wire                io_axi_25_aw_valid            ;
wire      [32:0]    io_axi_25_aw_bits_addr        ;
wire      [1:0]     io_axi_25_aw_bits_burst       ;
wire      [3:0]     io_axi_25_aw_bits_cache       ;
wire      [5:0]     io_axi_25_aw_bits_id          ;
wire      [3:0]     io_axi_25_aw_bits_len         ;
wire                io_axi_25_aw_bits_lock        ;
wire      [2:0]     io_axi_25_aw_bits_prot        ;
wire      [3:0]     io_axi_25_aw_bits_qos         ;
wire      [3:0]     io_axi_25_aw_bits_region      ;
wire      [2:0]     io_axi_25_aw_bits_size        ;
reg                 io_axi_25_ar_ready            =0;
wire                io_axi_25_ar_valid            ;
wire      [32:0]    io_axi_25_ar_bits_addr        ;
wire      [1:0]     io_axi_25_ar_bits_burst       ;
wire      [3:0]     io_axi_25_ar_bits_cache       ;
wire      [5:0]     io_axi_25_ar_bits_id          ;
wire      [3:0]     io_axi_25_ar_bits_len         ;
wire                io_axi_25_ar_bits_lock        ;
wire      [2:0]     io_axi_25_ar_bits_prot        ;
wire      [3:0]     io_axi_25_ar_bits_qos         ;
wire      [3:0]     io_axi_25_ar_bits_region      ;
wire      [2:0]     io_axi_25_ar_bits_size        ;
reg                 io_axi_25_w_ready             =0;
wire                io_axi_25_w_valid             ;
wire      [255:0]   io_axi_25_w_bits_data         ;
wire                io_axi_25_w_bits_last         ;
wire      [31:0]    io_axi_25_w_bits_strb         ;
wire                io_axi_25_r_ready             ;
reg                 io_axi_25_r_valid             =0;
reg       [255:0]   io_axi_25_r_bits_data         =0;
reg                 io_axi_25_r_bits_last         =0;
reg       [1:0]     io_axi_25_r_bits_resp         =0;
reg       [5:0]     io_axi_25_r_bits_id           =0;
wire                io_axi_25_b_ready             ;
reg                 io_axi_25_b_valid             =0;
reg       [5:0]     io_axi_25_b_bits_id           =0;
reg       [1:0]     io_axi_25_b_bits_resp         =0;
reg                 io_axi_26_aw_ready            =0;
wire                io_axi_26_aw_valid            ;
wire      [32:0]    io_axi_26_aw_bits_addr        ;
wire      [1:0]     io_axi_26_aw_bits_burst       ;
wire      [3:0]     io_axi_26_aw_bits_cache       ;
wire      [5:0]     io_axi_26_aw_bits_id          ;
wire      [3:0]     io_axi_26_aw_bits_len         ;
wire                io_axi_26_aw_bits_lock        ;
wire      [2:0]     io_axi_26_aw_bits_prot        ;
wire      [3:0]     io_axi_26_aw_bits_qos         ;
wire      [3:0]     io_axi_26_aw_bits_region      ;
wire      [2:0]     io_axi_26_aw_bits_size        ;
reg                 io_axi_26_ar_ready            =0;
wire                io_axi_26_ar_valid            ;
wire      [32:0]    io_axi_26_ar_bits_addr        ;
wire      [1:0]     io_axi_26_ar_bits_burst       ;
wire      [3:0]     io_axi_26_ar_bits_cache       ;
wire      [5:0]     io_axi_26_ar_bits_id          ;
wire      [3:0]     io_axi_26_ar_bits_len         ;
wire                io_axi_26_ar_bits_lock        ;
wire      [2:0]     io_axi_26_ar_bits_prot        ;
wire      [3:0]     io_axi_26_ar_bits_qos         ;
wire      [3:0]     io_axi_26_ar_bits_region      ;
wire      [2:0]     io_axi_26_ar_bits_size        ;
reg                 io_axi_26_w_ready             =0;
wire                io_axi_26_w_valid             ;
wire      [255:0]   io_axi_26_w_bits_data         ;
wire                io_axi_26_w_bits_last         ;
wire      [31:0]    io_axi_26_w_bits_strb         ;
wire                io_axi_26_r_ready             ;
reg                 io_axi_26_r_valid             =0;
reg       [255:0]   io_axi_26_r_bits_data         =0;
reg                 io_axi_26_r_bits_last         =0;
reg       [1:0]     io_axi_26_r_bits_resp         =0;
reg       [5:0]     io_axi_26_r_bits_id           =0;
wire                io_axi_26_b_ready             ;
reg                 io_axi_26_b_valid             =0;
reg       [5:0]     io_axi_26_b_bits_id           =0;
reg       [1:0]     io_axi_26_b_bits_resp         =0;
reg                 io_axi_27_aw_ready            =0;
wire                io_axi_27_aw_valid            ;
wire      [32:0]    io_axi_27_aw_bits_addr        ;
wire      [1:0]     io_axi_27_aw_bits_burst       ;
wire      [3:0]     io_axi_27_aw_bits_cache       ;
wire      [5:0]     io_axi_27_aw_bits_id          ;
wire      [3:0]     io_axi_27_aw_bits_len         ;
wire                io_axi_27_aw_bits_lock        ;
wire      [2:0]     io_axi_27_aw_bits_prot        ;
wire      [3:0]     io_axi_27_aw_bits_qos         ;
wire      [3:0]     io_axi_27_aw_bits_region      ;
wire      [2:0]     io_axi_27_aw_bits_size        ;
reg                 io_axi_27_ar_ready            =0;
wire                io_axi_27_ar_valid            ;
wire      [32:0]    io_axi_27_ar_bits_addr        ;
wire      [1:0]     io_axi_27_ar_bits_burst       ;
wire      [3:0]     io_axi_27_ar_bits_cache       ;
wire      [5:0]     io_axi_27_ar_bits_id          ;
wire      [3:0]     io_axi_27_ar_bits_len         ;
wire                io_axi_27_ar_bits_lock        ;
wire      [2:0]     io_axi_27_ar_bits_prot        ;
wire      [3:0]     io_axi_27_ar_bits_qos         ;
wire      [3:0]     io_axi_27_ar_bits_region      ;
wire      [2:0]     io_axi_27_ar_bits_size        ;
reg                 io_axi_27_w_ready             =0;
wire                io_axi_27_w_valid             ;
wire      [255:0]   io_axi_27_w_bits_data         ;
wire                io_axi_27_w_bits_last         ;
wire      [31:0]    io_axi_27_w_bits_strb         ;
wire                io_axi_27_r_ready             ;
reg                 io_axi_27_r_valid             =0;
reg       [255:0]   io_axi_27_r_bits_data         =0;
reg                 io_axi_27_r_bits_last         =0;
reg       [1:0]     io_axi_27_r_bits_resp         =0;
reg       [5:0]     io_axi_27_r_bits_id           =0;
wire                io_axi_27_b_ready             ;
reg                 io_axi_27_b_valid             =0;
reg       [5:0]     io_axi_27_b_bits_id           =0;
reg       [1:0]     io_axi_27_b_bits_resp         =0;
reg                 io_axi_28_aw_ready            =0;
wire                io_axi_28_aw_valid            ;
wire      [32:0]    io_axi_28_aw_bits_addr        ;
wire      [1:0]     io_axi_28_aw_bits_burst       ;
wire      [3:0]     io_axi_28_aw_bits_cache       ;
wire      [5:0]     io_axi_28_aw_bits_id          ;
wire      [3:0]     io_axi_28_aw_bits_len         ;
wire                io_axi_28_aw_bits_lock        ;
wire      [2:0]     io_axi_28_aw_bits_prot        ;
wire      [3:0]     io_axi_28_aw_bits_qos         ;
wire      [3:0]     io_axi_28_aw_bits_region      ;
wire      [2:0]     io_axi_28_aw_bits_size        ;
reg                 io_axi_28_ar_ready            =0;
wire                io_axi_28_ar_valid            ;
wire      [32:0]    io_axi_28_ar_bits_addr        ;
wire      [1:0]     io_axi_28_ar_bits_burst       ;
wire      [3:0]     io_axi_28_ar_bits_cache       ;
wire      [5:0]     io_axi_28_ar_bits_id          ;
wire      [3:0]     io_axi_28_ar_bits_len         ;
wire                io_axi_28_ar_bits_lock        ;
wire      [2:0]     io_axi_28_ar_bits_prot        ;
wire      [3:0]     io_axi_28_ar_bits_qos         ;
wire      [3:0]     io_axi_28_ar_bits_region      ;
wire      [2:0]     io_axi_28_ar_bits_size        ;
reg                 io_axi_28_w_ready             =0;
wire                io_axi_28_w_valid             ;
wire      [255:0]   io_axi_28_w_bits_data         ;
wire                io_axi_28_w_bits_last         ;
wire      [31:0]    io_axi_28_w_bits_strb         ;
wire                io_axi_28_r_ready             ;
reg                 io_axi_28_r_valid             =0;
reg       [255:0]   io_axi_28_r_bits_data         =0;
reg                 io_axi_28_r_bits_last         =0;
reg       [1:0]     io_axi_28_r_bits_resp         =0;
reg       [5:0]     io_axi_28_r_bits_id           =0;
wire                io_axi_28_b_ready             ;
reg                 io_axi_28_b_valid             =0;
reg       [5:0]     io_axi_28_b_bits_id           =0;
reg       [1:0]     io_axi_28_b_bits_resp         =0;
reg                 io_axi_29_aw_ready            =0;
wire                io_axi_29_aw_valid            ;
wire      [32:0]    io_axi_29_aw_bits_addr        ;
wire      [1:0]     io_axi_29_aw_bits_burst       ;
wire      [3:0]     io_axi_29_aw_bits_cache       ;
wire      [5:0]     io_axi_29_aw_bits_id          ;
wire      [3:0]     io_axi_29_aw_bits_len         ;
wire                io_axi_29_aw_bits_lock        ;
wire      [2:0]     io_axi_29_aw_bits_prot        ;
wire      [3:0]     io_axi_29_aw_bits_qos         ;
wire      [3:0]     io_axi_29_aw_bits_region      ;
wire      [2:0]     io_axi_29_aw_bits_size        ;
reg                 io_axi_29_ar_ready            =0;
wire                io_axi_29_ar_valid            ;
wire      [32:0]    io_axi_29_ar_bits_addr        ;
wire      [1:0]     io_axi_29_ar_bits_burst       ;
wire      [3:0]     io_axi_29_ar_bits_cache       ;
wire      [5:0]     io_axi_29_ar_bits_id          ;
wire      [3:0]     io_axi_29_ar_bits_len         ;
wire                io_axi_29_ar_bits_lock        ;
wire      [2:0]     io_axi_29_ar_bits_prot        ;
wire      [3:0]     io_axi_29_ar_bits_qos         ;
wire      [3:0]     io_axi_29_ar_bits_region      ;
wire      [2:0]     io_axi_29_ar_bits_size        ;
reg                 io_axi_29_w_ready             =0;
wire                io_axi_29_w_valid             ;
wire      [255:0]   io_axi_29_w_bits_data         ;
wire                io_axi_29_w_bits_last         ;
wire      [31:0]    io_axi_29_w_bits_strb         ;
wire                io_axi_29_r_ready             ;
reg                 io_axi_29_r_valid             =0;
reg       [255:0]   io_axi_29_r_bits_data         =0;
reg                 io_axi_29_r_bits_last         =0;
reg       [1:0]     io_axi_29_r_bits_resp         =0;
reg       [5:0]     io_axi_29_r_bits_id           =0;
wire                io_axi_29_b_ready             ;
reg                 io_axi_29_b_valid             =0;
reg       [5:0]     io_axi_29_b_bits_id           =0;
reg       [1:0]     io_axi_29_b_bits_resp         =0;
reg                 io_axi_30_aw_ready            =0;
wire                io_axi_30_aw_valid            ;
wire      [32:0]    io_axi_30_aw_bits_addr        ;
wire      [1:0]     io_axi_30_aw_bits_burst       ;
wire      [3:0]     io_axi_30_aw_bits_cache       ;
wire      [5:0]     io_axi_30_aw_bits_id          ;
wire      [3:0]     io_axi_30_aw_bits_len         ;
wire                io_axi_30_aw_bits_lock        ;
wire      [2:0]     io_axi_30_aw_bits_prot        ;
wire      [3:0]     io_axi_30_aw_bits_qos         ;
wire      [3:0]     io_axi_30_aw_bits_region      ;
wire      [2:0]     io_axi_30_aw_bits_size        ;
reg                 io_axi_30_ar_ready            =0;
wire                io_axi_30_ar_valid            ;
wire      [32:0]    io_axi_30_ar_bits_addr        ;
wire      [1:0]     io_axi_30_ar_bits_burst       ;
wire      [3:0]     io_axi_30_ar_bits_cache       ;
wire      [5:0]     io_axi_30_ar_bits_id          ;
wire      [3:0]     io_axi_30_ar_bits_len         ;
wire                io_axi_30_ar_bits_lock        ;
wire      [2:0]     io_axi_30_ar_bits_prot        ;
wire      [3:0]     io_axi_30_ar_bits_qos         ;
wire      [3:0]     io_axi_30_ar_bits_region      ;
wire      [2:0]     io_axi_30_ar_bits_size        ;
reg                 io_axi_30_w_ready             =0;
wire                io_axi_30_w_valid             ;
wire      [255:0]   io_axi_30_w_bits_data         ;
wire                io_axi_30_w_bits_last         ;
wire      [31:0]    io_axi_30_w_bits_strb         ;
wire                io_axi_30_r_ready             ;
reg                 io_axi_30_r_valid             =0;
reg       [255:0]   io_axi_30_r_bits_data         =0;
reg                 io_axi_30_r_bits_last         =0;
reg       [1:0]     io_axi_30_r_bits_resp         =0;
reg       [5:0]     io_axi_30_r_bits_id           =0;
wire                io_axi_30_b_ready             ;
reg                 io_axi_30_b_valid             =0;
reg       [5:0]     io_axi_30_b_bits_id           =0;
reg       [1:0]     io_axi_30_b_bits_resp         =0;
reg                 io_axi_31_aw_ready            =0;
wire                io_axi_31_aw_valid            ;
wire      [32:0]    io_axi_31_aw_bits_addr        ;
wire      [1:0]     io_axi_31_aw_bits_burst       ;
wire      [3:0]     io_axi_31_aw_bits_cache       ;
wire      [5:0]     io_axi_31_aw_bits_id          ;
wire      [3:0]     io_axi_31_aw_bits_len         ;
wire                io_axi_31_aw_bits_lock        ;
wire      [2:0]     io_axi_31_aw_bits_prot        ;
wire      [3:0]     io_axi_31_aw_bits_qos         ;
wire      [3:0]     io_axi_31_aw_bits_region      ;
wire      [2:0]     io_axi_31_aw_bits_size        ;
reg                 io_axi_31_ar_ready            =0;
wire                io_axi_31_ar_valid            ;
wire      [32:0]    io_axi_31_ar_bits_addr        ;
wire      [1:0]     io_axi_31_ar_bits_burst       ;
wire      [3:0]     io_axi_31_ar_bits_cache       ;
wire      [5:0]     io_axi_31_ar_bits_id          ;
wire      [3:0]     io_axi_31_ar_bits_len         ;
wire                io_axi_31_ar_bits_lock        ;
wire      [2:0]     io_axi_31_ar_bits_prot        ;
wire      [3:0]     io_axi_31_ar_bits_qos         ;
wire      [3:0]     io_axi_31_ar_bits_region      ;
wire      [2:0]     io_axi_31_ar_bits_size        ;
reg                 io_axi_31_w_ready             =0;
wire                io_axi_31_w_valid             ;
wire      [255:0]   io_axi_31_w_bits_data         ;
wire                io_axi_31_w_bits_last         ;
wire      [31:0]    io_axi_31_w_bits_strb         ;
wire                io_axi_31_r_ready             ;
reg                 io_axi_31_r_valid             =0;
reg       [255:0]   io_axi_31_r_bits_data         =0;
reg                 io_axi_31_r_bits_last         =0;
reg       [1:0]     io_axi_31_r_bits_resp         =0;
reg       [5:0]     io_axi_31_r_bits_id           =0;
wire                io_axi_31_b_ready             ;
reg                 io_axi_31_b_valid             =0;
reg       [5:0]     io_axi_31_b_bits_id           =0;
reg       [1:0]     io_axi_31_b_bits_resp         =0;
reg                 io_start                      =0;
reg                 io_start_compress             =0;

OUT#(64)out_io_axi_0_aw(
        clock,
        reset,
        {io_axi_0_aw_bits_addr,io_axi_0_aw_bits_burst,io_axi_0_aw_bits_cache,io_axi_0_aw_bits_id,io_axi_0_aw_bits_len,io_axi_0_aw_bits_lock,io_axi_0_aw_bits_prot,io_axi_0_aw_bits_qos,io_axi_0_aw_bits_region,io_axi_0_aw_bits_size},
        io_axi_0_aw_valid,
        io_axi_0_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_0_ar(
        clock,
        reset,
        {io_axi_0_ar_bits_addr,io_axi_0_ar_bits_burst,io_axi_0_ar_bits_cache,io_axi_0_ar_bits_id,io_axi_0_ar_bits_len,io_axi_0_ar_bits_lock,io_axi_0_ar_bits_prot,io_axi_0_ar_bits_qos,io_axi_0_ar_bits_region,io_axi_0_ar_bits_size},
        io_axi_0_ar_valid,
        io_axi_0_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_0_w(
        clock,
        reset,
        {io_axi_0_w_bits_data,io_axi_0_w_bits_last,io_axi_0_w_bits_strb},
        io_axi_0_w_valid,
        io_axi_0_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_0_r(
        clock,
        reset,
        {io_axi_0_r_bits_data,io_axi_0_r_bits_last,io_axi_0_r_bits_resp,io_axi_0_r_bits_id},
        io_axi_0_r_valid,
        io_axi_0_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_0_b(
        clock,
        reset,
        {io_axi_0_b_bits_id,io_axi_0_b_bits_resp},
        io_axi_0_b_valid,
        io_axi_0_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_1_aw(
        clock,
        reset,
        {io_axi_1_aw_bits_addr,io_axi_1_aw_bits_burst,io_axi_1_aw_bits_cache,io_axi_1_aw_bits_id,io_axi_1_aw_bits_len,io_axi_1_aw_bits_lock,io_axi_1_aw_bits_prot,io_axi_1_aw_bits_qos,io_axi_1_aw_bits_region,io_axi_1_aw_bits_size},
        io_axi_1_aw_valid,
        io_axi_1_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_1_ar(
        clock,
        reset,
        {io_axi_1_ar_bits_addr,io_axi_1_ar_bits_burst,io_axi_1_ar_bits_cache,io_axi_1_ar_bits_id,io_axi_1_ar_bits_len,io_axi_1_ar_bits_lock,io_axi_1_ar_bits_prot,io_axi_1_ar_bits_qos,io_axi_1_ar_bits_region,io_axi_1_ar_bits_size},
        io_axi_1_ar_valid,
        io_axi_1_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_1_w(
        clock,
        reset,
        {io_axi_1_w_bits_data,io_axi_1_w_bits_last,io_axi_1_w_bits_strb},
        io_axi_1_w_valid,
        io_axi_1_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_1_r(
        clock,
        reset,
        {io_axi_1_r_bits_data,io_axi_1_r_bits_last,io_axi_1_r_bits_resp,io_axi_1_r_bits_id},
        io_axi_1_r_valid,
        io_axi_1_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_1_b(
        clock,
        reset,
        {io_axi_1_b_bits_id,io_axi_1_b_bits_resp},
        io_axi_1_b_valid,
        io_axi_1_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_2_aw(
        clock,
        reset,
        {io_axi_2_aw_bits_addr,io_axi_2_aw_bits_burst,io_axi_2_aw_bits_cache,io_axi_2_aw_bits_id,io_axi_2_aw_bits_len,io_axi_2_aw_bits_lock,io_axi_2_aw_bits_prot,io_axi_2_aw_bits_qos,io_axi_2_aw_bits_region,io_axi_2_aw_bits_size},
        io_axi_2_aw_valid,
        io_axi_2_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_2_ar(
        clock,
        reset,
        {io_axi_2_ar_bits_addr,io_axi_2_ar_bits_burst,io_axi_2_ar_bits_cache,io_axi_2_ar_bits_id,io_axi_2_ar_bits_len,io_axi_2_ar_bits_lock,io_axi_2_ar_bits_prot,io_axi_2_ar_bits_qos,io_axi_2_ar_bits_region,io_axi_2_ar_bits_size},
        io_axi_2_ar_valid,
        io_axi_2_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_2_w(
        clock,
        reset,
        {io_axi_2_w_bits_data,io_axi_2_w_bits_last,io_axi_2_w_bits_strb},
        io_axi_2_w_valid,
        io_axi_2_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_2_r(
        clock,
        reset,
        {io_axi_2_r_bits_data,io_axi_2_r_bits_last,io_axi_2_r_bits_resp,io_axi_2_r_bits_id},
        io_axi_2_r_valid,
        io_axi_2_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_2_b(
        clock,
        reset,
        {io_axi_2_b_bits_id,io_axi_2_b_bits_resp},
        io_axi_2_b_valid,
        io_axi_2_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_3_aw(
        clock,
        reset,
        {io_axi_3_aw_bits_addr,io_axi_3_aw_bits_burst,io_axi_3_aw_bits_cache,io_axi_3_aw_bits_id,io_axi_3_aw_bits_len,io_axi_3_aw_bits_lock,io_axi_3_aw_bits_prot,io_axi_3_aw_bits_qos,io_axi_3_aw_bits_region,io_axi_3_aw_bits_size},
        io_axi_3_aw_valid,
        io_axi_3_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_3_ar(
        clock,
        reset,
        {io_axi_3_ar_bits_addr,io_axi_3_ar_bits_burst,io_axi_3_ar_bits_cache,io_axi_3_ar_bits_id,io_axi_3_ar_bits_len,io_axi_3_ar_bits_lock,io_axi_3_ar_bits_prot,io_axi_3_ar_bits_qos,io_axi_3_ar_bits_region,io_axi_3_ar_bits_size},
        io_axi_3_ar_valid,
        io_axi_3_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_3_w(
        clock,
        reset,
        {io_axi_3_w_bits_data,io_axi_3_w_bits_last,io_axi_3_w_bits_strb},
        io_axi_3_w_valid,
        io_axi_3_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_3_r(
        clock,
        reset,
        {io_axi_3_r_bits_data,io_axi_3_r_bits_last,io_axi_3_r_bits_resp,io_axi_3_r_bits_id},
        io_axi_3_r_valid,
        io_axi_3_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_3_b(
        clock,
        reset,
        {io_axi_3_b_bits_id,io_axi_3_b_bits_resp},
        io_axi_3_b_valid,
        io_axi_3_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_4_aw(
        clock,
        reset,
        {io_axi_4_aw_bits_addr,io_axi_4_aw_bits_burst,io_axi_4_aw_bits_cache,io_axi_4_aw_bits_id,io_axi_4_aw_bits_len,io_axi_4_aw_bits_lock,io_axi_4_aw_bits_prot,io_axi_4_aw_bits_qos,io_axi_4_aw_bits_region,io_axi_4_aw_bits_size},
        io_axi_4_aw_valid,
        io_axi_4_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_4_ar(
        clock,
        reset,
        {io_axi_4_ar_bits_addr,io_axi_4_ar_bits_burst,io_axi_4_ar_bits_cache,io_axi_4_ar_bits_id,io_axi_4_ar_bits_len,io_axi_4_ar_bits_lock,io_axi_4_ar_bits_prot,io_axi_4_ar_bits_qos,io_axi_4_ar_bits_region,io_axi_4_ar_bits_size},
        io_axi_4_ar_valid,
        io_axi_4_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_4_w(
        clock,
        reset,
        {io_axi_4_w_bits_data,io_axi_4_w_bits_last,io_axi_4_w_bits_strb},
        io_axi_4_w_valid,
        io_axi_4_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_4_r(
        clock,
        reset,
        {io_axi_4_r_bits_data,io_axi_4_r_bits_last,io_axi_4_r_bits_resp,io_axi_4_r_bits_id},
        io_axi_4_r_valid,
        io_axi_4_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_4_b(
        clock,
        reset,
        {io_axi_4_b_bits_id,io_axi_4_b_bits_resp},
        io_axi_4_b_valid,
        io_axi_4_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_5_aw(
        clock,
        reset,
        {io_axi_5_aw_bits_addr,io_axi_5_aw_bits_burst,io_axi_5_aw_bits_cache,io_axi_5_aw_bits_id,io_axi_5_aw_bits_len,io_axi_5_aw_bits_lock,io_axi_5_aw_bits_prot,io_axi_5_aw_bits_qos,io_axi_5_aw_bits_region,io_axi_5_aw_bits_size},
        io_axi_5_aw_valid,
        io_axi_5_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_5_ar(
        clock,
        reset,
        {io_axi_5_ar_bits_addr,io_axi_5_ar_bits_burst,io_axi_5_ar_bits_cache,io_axi_5_ar_bits_id,io_axi_5_ar_bits_len,io_axi_5_ar_bits_lock,io_axi_5_ar_bits_prot,io_axi_5_ar_bits_qos,io_axi_5_ar_bits_region,io_axi_5_ar_bits_size},
        io_axi_5_ar_valid,
        io_axi_5_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_5_w(
        clock,
        reset,
        {io_axi_5_w_bits_data,io_axi_5_w_bits_last,io_axi_5_w_bits_strb},
        io_axi_5_w_valid,
        io_axi_5_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_5_r(
        clock,
        reset,
        {io_axi_5_r_bits_data,io_axi_5_r_bits_last,io_axi_5_r_bits_resp,io_axi_5_r_bits_id},
        io_axi_5_r_valid,
        io_axi_5_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_5_b(
        clock,
        reset,
        {io_axi_5_b_bits_id,io_axi_5_b_bits_resp},
        io_axi_5_b_valid,
        io_axi_5_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_6_aw(
        clock,
        reset,
        {io_axi_6_aw_bits_addr,io_axi_6_aw_bits_burst,io_axi_6_aw_bits_cache,io_axi_6_aw_bits_id,io_axi_6_aw_bits_len,io_axi_6_aw_bits_lock,io_axi_6_aw_bits_prot,io_axi_6_aw_bits_qos,io_axi_6_aw_bits_region,io_axi_6_aw_bits_size},
        io_axi_6_aw_valid,
        io_axi_6_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_6_ar(
        clock,
        reset,
        {io_axi_6_ar_bits_addr,io_axi_6_ar_bits_burst,io_axi_6_ar_bits_cache,io_axi_6_ar_bits_id,io_axi_6_ar_bits_len,io_axi_6_ar_bits_lock,io_axi_6_ar_bits_prot,io_axi_6_ar_bits_qos,io_axi_6_ar_bits_region,io_axi_6_ar_bits_size},
        io_axi_6_ar_valid,
        io_axi_6_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_6_w(
        clock,
        reset,
        {io_axi_6_w_bits_data,io_axi_6_w_bits_last,io_axi_6_w_bits_strb},
        io_axi_6_w_valid,
        io_axi_6_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_6_r(
        clock,
        reset,
        {io_axi_6_r_bits_data,io_axi_6_r_bits_last,io_axi_6_r_bits_resp,io_axi_6_r_bits_id},
        io_axi_6_r_valid,
        io_axi_6_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_6_b(
        clock,
        reset,
        {io_axi_6_b_bits_id,io_axi_6_b_bits_resp},
        io_axi_6_b_valid,
        io_axi_6_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_7_aw(
        clock,
        reset,
        {io_axi_7_aw_bits_addr,io_axi_7_aw_bits_burst,io_axi_7_aw_bits_cache,io_axi_7_aw_bits_id,io_axi_7_aw_bits_len,io_axi_7_aw_bits_lock,io_axi_7_aw_bits_prot,io_axi_7_aw_bits_qos,io_axi_7_aw_bits_region,io_axi_7_aw_bits_size},
        io_axi_7_aw_valid,
        io_axi_7_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_7_ar(
        clock,
        reset,
        {io_axi_7_ar_bits_addr,io_axi_7_ar_bits_burst,io_axi_7_ar_bits_cache,io_axi_7_ar_bits_id,io_axi_7_ar_bits_len,io_axi_7_ar_bits_lock,io_axi_7_ar_bits_prot,io_axi_7_ar_bits_qos,io_axi_7_ar_bits_region,io_axi_7_ar_bits_size},
        io_axi_7_ar_valid,
        io_axi_7_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_7_w(
        clock,
        reset,
        {io_axi_7_w_bits_data,io_axi_7_w_bits_last,io_axi_7_w_bits_strb},
        io_axi_7_w_valid,
        io_axi_7_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_7_r(
        clock,
        reset,
        {io_axi_7_r_bits_data,io_axi_7_r_bits_last,io_axi_7_r_bits_resp,io_axi_7_r_bits_id},
        io_axi_7_r_valid,
        io_axi_7_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_7_b(
        clock,
        reset,
        {io_axi_7_b_bits_id,io_axi_7_b_bits_resp},
        io_axi_7_b_valid,
        io_axi_7_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_8_aw(
        clock,
        reset,
        {io_axi_8_aw_bits_addr,io_axi_8_aw_bits_burst,io_axi_8_aw_bits_cache,io_axi_8_aw_bits_id,io_axi_8_aw_bits_len,io_axi_8_aw_bits_lock,io_axi_8_aw_bits_prot,io_axi_8_aw_bits_qos,io_axi_8_aw_bits_region,io_axi_8_aw_bits_size},
        io_axi_8_aw_valid,
        io_axi_8_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_8_ar(
        clock,
        reset,
        {io_axi_8_ar_bits_addr,io_axi_8_ar_bits_burst,io_axi_8_ar_bits_cache,io_axi_8_ar_bits_id,io_axi_8_ar_bits_len,io_axi_8_ar_bits_lock,io_axi_8_ar_bits_prot,io_axi_8_ar_bits_qos,io_axi_8_ar_bits_region,io_axi_8_ar_bits_size},
        io_axi_8_ar_valid,
        io_axi_8_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_8_w(
        clock,
        reset,
        {io_axi_8_w_bits_data,io_axi_8_w_bits_last,io_axi_8_w_bits_strb},
        io_axi_8_w_valid,
        io_axi_8_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_8_r(
        clock,
        reset,
        {io_axi_8_r_bits_data,io_axi_8_r_bits_last,io_axi_8_r_bits_resp,io_axi_8_r_bits_id},
        io_axi_8_r_valid,
        io_axi_8_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_8_b(
        clock,
        reset,
        {io_axi_8_b_bits_id,io_axi_8_b_bits_resp},
        io_axi_8_b_valid,
        io_axi_8_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_9_aw(
        clock,
        reset,
        {io_axi_9_aw_bits_addr,io_axi_9_aw_bits_burst,io_axi_9_aw_bits_cache,io_axi_9_aw_bits_id,io_axi_9_aw_bits_len,io_axi_9_aw_bits_lock,io_axi_9_aw_bits_prot,io_axi_9_aw_bits_qos,io_axi_9_aw_bits_region,io_axi_9_aw_bits_size},
        io_axi_9_aw_valid,
        io_axi_9_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_9_ar(
        clock,
        reset,
        {io_axi_9_ar_bits_addr,io_axi_9_ar_bits_burst,io_axi_9_ar_bits_cache,io_axi_9_ar_bits_id,io_axi_9_ar_bits_len,io_axi_9_ar_bits_lock,io_axi_9_ar_bits_prot,io_axi_9_ar_bits_qos,io_axi_9_ar_bits_region,io_axi_9_ar_bits_size},
        io_axi_9_ar_valid,
        io_axi_9_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_9_w(
        clock,
        reset,
        {io_axi_9_w_bits_data,io_axi_9_w_bits_last,io_axi_9_w_bits_strb},
        io_axi_9_w_valid,
        io_axi_9_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_9_r(
        clock,
        reset,
        {io_axi_9_r_bits_data,io_axi_9_r_bits_last,io_axi_9_r_bits_resp,io_axi_9_r_bits_id},
        io_axi_9_r_valid,
        io_axi_9_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_9_b(
        clock,
        reset,
        {io_axi_9_b_bits_id,io_axi_9_b_bits_resp},
        io_axi_9_b_valid,
        io_axi_9_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_10_aw(
        clock,
        reset,
        {io_axi_10_aw_bits_addr,io_axi_10_aw_bits_burst,io_axi_10_aw_bits_cache,io_axi_10_aw_bits_id,io_axi_10_aw_bits_len,io_axi_10_aw_bits_lock,io_axi_10_aw_bits_prot,io_axi_10_aw_bits_qos,io_axi_10_aw_bits_region,io_axi_10_aw_bits_size},
        io_axi_10_aw_valid,
        io_axi_10_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_10_ar(
        clock,
        reset,
        {io_axi_10_ar_bits_addr,io_axi_10_ar_bits_burst,io_axi_10_ar_bits_cache,io_axi_10_ar_bits_id,io_axi_10_ar_bits_len,io_axi_10_ar_bits_lock,io_axi_10_ar_bits_prot,io_axi_10_ar_bits_qos,io_axi_10_ar_bits_region,io_axi_10_ar_bits_size},
        io_axi_10_ar_valid,
        io_axi_10_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_10_w(
        clock,
        reset,
        {io_axi_10_w_bits_data,io_axi_10_w_bits_last,io_axi_10_w_bits_strb},
        io_axi_10_w_valid,
        io_axi_10_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_10_r(
        clock,
        reset,
        {io_axi_10_r_bits_data,io_axi_10_r_bits_last,io_axi_10_r_bits_resp,io_axi_10_r_bits_id},
        io_axi_10_r_valid,
        io_axi_10_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_10_b(
        clock,
        reset,
        {io_axi_10_b_bits_id,io_axi_10_b_bits_resp},
        io_axi_10_b_valid,
        io_axi_10_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_11_aw(
        clock,
        reset,
        {io_axi_11_aw_bits_addr,io_axi_11_aw_bits_burst,io_axi_11_aw_bits_cache,io_axi_11_aw_bits_id,io_axi_11_aw_bits_len,io_axi_11_aw_bits_lock,io_axi_11_aw_bits_prot,io_axi_11_aw_bits_qos,io_axi_11_aw_bits_region,io_axi_11_aw_bits_size},
        io_axi_11_aw_valid,
        io_axi_11_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_11_ar(
        clock,
        reset,
        {io_axi_11_ar_bits_addr,io_axi_11_ar_bits_burst,io_axi_11_ar_bits_cache,io_axi_11_ar_bits_id,io_axi_11_ar_bits_len,io_axi_11_ar_bits_lock,io_axi_11_ar_bits_prot,io_axi_11_ar_bits_qos,io_axi_11_ar_bits_region,io_axi_11_ar_bits_size},
        io_axi_11_ar_valid,
        io_axi_11_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_11_w(
        clock,
        reset,
        {io_axi_11_w_bits_data,io_axi_11_w_bits_last,io_axi_11_w_bits_strb},
        io_axi_11_w_valid,
        io_axi_11_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_11_r(
        clock,
        reset,
        {io_axi_11_r_bits_data,io_axi_11_r_bits_last,io_axi_11_r_bits_resp,io_axi_11_r_bits_id},
        io_axi_11_r_valid,
        io_axi_11_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_11_b(
        clock,
        reset,
        {io_axi_11_b_bits_id,io_axi_11_b_bits_resp},
        io_axi_11_b_valid,
        io_axi_11_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_12_aw(
        clock,
        reset,
        {io_axi_12_aw_bits_addr,io_axi_12_aw_bits_burst,io_axi_12_aw_bits_cache,io_axi_12_aw_bits_id,io_axi_12_aw_bits_len,io_axi_12_aw_bits_lock,io_axi_12_aw_bits_prot,io_axi_12_aw_bits_qos,io_axi_12_aw_bits_region,io_axi_12_aw_bits_size},
        io_axi_12_aw_valid,
        io_axi_12_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_12_ar(
        clock,
        reset,
        {io_axi_12_ar_bits_addr,io_axi_12_ar_bits_burst,io_axi_12_ar_bits_cache,io_axi_12_ar_bits_id,io_axi_12_ar_bits_len,io_axi_12_ar_bits_lock,io_axi_12_ar_bits_prot,io_axi_12_ar_bits_qos,io_axi_12_ar_bits_region,io_axi_12_ar_bits_size},
        io_axi_12_ar_valid,
        io_axi_12_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_12_w(
        clock,
        reset,
        {io_axi_12_w_bits_data,io_axi_12_w_bits_last,io_axi_12_w_bits_strb},
        io_axi_12_w_valid,
        io_axi_12_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_12_r(
        clock,
        reset,
        {io_axi_12_r_bits_data,io_axi_12_r_bits_last,io_axi_12_r_bits_resp,io_axi_12_r_bits_id},
        io_axi_12_r_valid,
        io_axi_12_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_12_b(
        clock,
        reset,
        {io_axi_12_b_bits_id,io_axi_12_b_bits_resp},
        io_axi_12_b_valid,
        io_axi_12_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_13_aw(
        clock,
        reset,
        {io_axi_13_aw_bits_addr,io_axi_13_aw_bits_burst,io_axi_13_aw_bits_cache,io_axi_13_aw_bits_id,io_axi_13_aw_bits_len,io_axi_13_aw_bits_lock,io_axi_13_aw_bits_prot,io_axi_13_aw_bits_qos,io_axi_13_aw_bits_region,io_axi_13_aw_bits_size},
        io_axi_13_aw_valid,
        io_axi_13_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_13_ar(
        clock,
        reset,
        {io_axi_13_ar_bits_addr,io_axi_13_ar_bits_burst,io_axi_13_ar_bits_cache,io_axi_13_ar_bits_id,io_axi_13_ar_bits_len,io_axi_13_ar_bits_lock,io_axi_13_ar_bits_prot,io_axi_13_ar_bits_qos,io_axi_13_ar_bits_region,io_axi_13_ar_bits_size},
        io_axi_13_ar_valid,
        io_axi_13_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_13_w(
        clock,
        reset,
        {io_axi_13_w_bits_data,io_axi_13_w_bits_last,io_axi_13_w_bits_strb},
        io_axi_13_w_valid,
        io_axi_13_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_13_r(
        clock,
        reset,
        {io_axi_13_r_bits_data,io_axi_13_r_bits_last,io_axi_13_r_bits_resp,io_axi_13_r_bits_id},
        io_axi_13_r_valid,
        io_axi_13_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_13_b(
        clock,
        reset,
        {io_axi_13_b_bits_id,io_axi_13_b_bits_resp},
        io_axi_13_b_valid,
        io_axi_13_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_14_aw(
        clock,
        reset,
        {io_axi_14_aw_bits_addr,io_axi_14_aw_bits_burst,io_axi_14_aw_bits_cache,io_axi_14_aw_bits_id,io_axi_14_aw_bits_len,io_axi_14_aw_bits_lock,io_axi_14_aw_bits_prot,io_axi_14_aw_bits_qos,io_axi_14_aw_bits_region,io_axi_14_aw_bits_size},
        io_axi_14_aw_valid,
        io_axi_14_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_14_ar(
        clock,
        reset,
        {io_axi_14_ar_bits_addr,io_axi_14_ar_bits_burst,io_axi_14_ar_bits_cache,io_axi_14_ar_bits_id,io_axi_14_ar_bits_len,io_axi_14_ar_bits_lock,io_axi_14_ar_bits_prot,io_axi_14_ar_bits_qos,io_axi_14_ar_bits_region,io_axi_14_ar_bits_size},
        io_axi_14_ar_valid,
        io_axi_14_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_14_w(
        clock,
        reset,
        {io_axi_14_w_bits_data,io_axi_14_w_bits_last,io_axi_14_w_bits_strb},
        io_axi_14_w_valid,
        io_axi_14_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_14_r(
        clock,
        reset,
        {io_axi_14_r_bits_data,io_axi_14_r_bits_last,io_axi_14_r_bits_resp,io_axi_14_r_bits_id},
        io_axi_14_r_valid,
        io_axi_14_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_14_b(
        clock,
        reset,
        {io_axi_14_b_bits_id,io_axi_14_b_bits_resp},
        io_axi_14_b_valid,
        io_axi_14_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_15_aw(
        clock,
        reset,
        {io_axi_15_aw_bits_addr,io_axi_15_aw_bits_burst,io_axi_15_aw_bits_cache,io_axi_15_aw_bits_id,io_axi_15_aw_bits_len,io_axi_15_aw_bits_lock,io_axi_15_aw_bits_prot,io_axi_15_aw_bits_qos,io_axi_15_aw_bits_region,io_axi_15_aw_bits_size},
        io_axi_15_aw_valid,
        io_axi_15_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_15_ar(
        clock,
        reset,
        {io_axi_15_ar_bits_addr,io_axi_15_ar_bits_burst,io_axi_15_ar_bits_cache,io_axi_15_ar_bits_id,io_axi_15_ar_bits_len,io_axi_15_ar_bits_lock,io_axi_15_ar_bits_prot,io_axi_15_ar_bits_qos,io_axi_15_ar_bits_region,io_axi_15_ar_bits_size},
        io_axi_15_ar_valid,
        io_axi_15_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_15_w(
        clock,
        reset,
        {io_axi_15_w_bits_data,io_axi_15_w_bits_last,io_axi_15_w_bits_strb},
        io_axi_15_w_valid,
        io_axi_15_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_15_r(
        clock,
        reset,
        {io_axi_15_r_bits_data,io_axi_15_r_bits_last,io_axi_15_r_bits_resp,io_axi_15_r_bits_id},
        io_axi_15_r_valid,
        io_axi_15_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_15_b(
        clock,
        reset,
        {io_axi_15_b_bits_id,io_axi_15_b_bits_resp},
        io_axi_15_b_valid,
        io_axi_15_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_16_aw(
        clock,
        reset,
        {io_axi_16_aw_bits_addr,io_axi_16_aw_bits_burst,io_axi_16_aw_bits_cache,io_axi_16_aw_bits_id,io_axi_16_aw_bits_len,io_axi_16_aw_bits_lock,io_axi_16_aw_bits_prot,io_axi_16_aw_bits_qos,io_axi_16_aw_bits_region,io_axi_16_aw_bits_size},
        io_axi_16_aw_valid,
        io_axi_16_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_16_ar(
        clock,
        reset,
        {io_axi_16_ar_bits_addr,io_axi_16_ar_bits_burst,io_axi_16_ar_bits_cache,io_axi_16_ar_bits_id,io_axi_16_ar_bits_len,io_axi_16_ar_bits_lock,io_axi_16_ar_bits_prot,io_axi_16_ar_bits_qos,io_axi_16_ar_bits_region,io_axi_16_ar_bits_size},
        io_axi_16_ar_valid,
        io_axi_16_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_16_w(
        clock,
        reset,
        {io_axi_16_w_bits_data,io_axi_16_w_bits_last,io_axi_16_w_bits_strb},
        io_axi_16_w_valid,
        io_axi_16_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_16_r(
        clock,
        reset,
        {io_axi_16_r_bits_data,io_axi_16_r_bits_last,io_axi_16_r_bits_resp,io_axi_16_r_bits_id},
        io_axi_16_r_valid,
        io_axi_16_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_16_b(
        clock,
        reset,
        {io_axi_16_b_bits_id,io_axi_16_b_bits_resp},
        io_axi_16_b_valid,
        io_axi_16_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_17_aw(
        clock,
        reset,
        {io_axi_17_aw_bits_addr,io_axi_17_aw_bits_burst,io_axi_17_aw_bits_cache,io_axi_17_aw_bits_id,io_axi_17_aw_bits_len,io_axi_17_aw_bits_lock,io_axi_17_aw_bits_prot,io_axi_17_aw_bits_qos,io_axi_17_aw_bits_region,io_axi_17_aw_bits_size},
        io_axi_17_aw_valid,
        io_axi_17_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_17_ar(
        clock,
        reset,
        {io_axi_17_ar_bits_addr,io_axi_17_ar_bits_burst,io_axi_17_ar_bits_cache,io_axi_17_ar_bits_id,io_axi_17_ar_bits_len,io_axi_17_ar_bits_lock,io_axi_17_ar_bits_prot,io_axi_17_ar_bits_qos,io_axi_17_ar_bits_region,io_axi_17_ar_bits_size},
        io_axi_17_ar_valid,
        io_axi_17_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_17_w(
        clock,
        reset,
        {io_axi_17_w_bits_data,io_axi_17_w_bits_last,io_axi_17_w_bits_strb},
        io_axi_17_w_valid,
        io_axi_17_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_17_r(
        clock,
        reset,
        {io_axi_17_r_bits_data,io_axi_17_r_bits_last,io_axi_17_r_bits_resp,io_axi_17_r_bits_id},
        io_axi_17_r_valid,
        io_axi_17_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_17_b(
        clock,
        reset,
        {io_axi_17_b_bits_id,io_axi_17_b_bits_resp},
        io_axi_17_b_valid,
        io_axi_17_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_18_aw(
        clock,
        reset,
        {io_axi_18_aw_bits_addr,io_axi_18_aw_bits_burst,io_axi_18_aw_bits_cache,io_axi_18_aw_bits_id,io_axi_18_aw_bits_len,io_axi_18_aw_bits_lock,io_axi_18_aw_bits_prot,io_axi_18_aw_bits_qos,io_axi_18_aw_bits_region,io_axi_18_aw_bits_size},
        io_axi_18_aw_valid,
        io_axi_18_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_18_ar(
        clock,
        reset,
        {io_axi_18_ar_bits_addr,io_axi_18_ar_bits_burst,io_axi_18_ar_bits_cache,io_axi_18_ar_bits_id,io_axi_18_ar_bits_len,io_axi_18_ar_bits_lock,io_axi_18_ar_bits_prot,io_axi_18_ar_bits_qos,io_axi_18_ar_bits_region,io_axi_18_ar_bits_size},
        io_axi_18_ar_valid,
        io_axi_18_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_18_w(
        clock,
        reset,
        {io_axi_18_w_bits_data,io_axi_18_w_bits_last,io_axi_18_w_bits_strb},
        io_axi_18_w_valid,
        io_axi_18_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_18_r(
        clock,
        reset,
        {io_axi_18_r_bits_data,io_axi_18_r_bits_last,io_axi_18_r_bits_resp,io_axi_18_r_bits_id},
        io_axi_18_r_valid,
        io_axi_18_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_18_b(
        clock,
        reset,
        {io_axi_18_b_bits_id,io_axi_18_b_bits_resp},
        io_axi_18_b_valid,
        io_axi_18_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_19_aw(
        clock,
        reset,
        {io_axi_19_aw_bits_addr,io_axi_19_aw_bits_burst,io_axi_19_aw_bits_cache,io_axi_19_aw_bits_id,io_axi_19_aw_bits_len,io_axi_19_aw_bits_lock,io_axi_19_aw_bits_prot,io_axi_19_aw_bits_qos,io_axi_19_aw_bits_region,io_axi_19_aw_bits_size},
        io_axi_19_aw_valid,
        io_axi_19_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_19_ar(
        clock,
        reset,
        {io_axi_19_ar_bits_addr,io_axi_19_ar_bits_burst,io_axi_19_ar_bits_cache,io_axi_19_ar_bits_id,io_axi_19_ar_bits_len,io_axi_19_ar_bits_lock,io_axi_19_ar_bits_prot,io_axi_19_ar_bits_qos,io_axi_19_ar_bits_region,io_axi_19_ar_bits_size},
        io_axi_19_ar_valid,
        io_axi_19_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_19_w(
        clock,
        reset,
        {io_axi_19_w_bits_data,io_axi_19_w_bits_last,io_axi_19_w_bits_strb},
        io_axi_19_w_valid,
        io_axi_19_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_19_r(
        clock,
        reset,
        {io_axi_19_r_bits_data,io_axi_19_r_bits_last,io_axi_19_r_bits_resp,io_axi_19_r_bits_id},
        io_axi_19_r_valid,
        io_axi_19_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_19_b(
        clock,
        reset,
        {io_axi_19_b_bits_id,io_axi_19_b_bits_resp},
        io_axi_19_b_valid,
        io_axi_19_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_20_aw(
        clock,
        reset,
        {io_axi_20_aw_bits_addr,io_axi_20_aw_bits_burst,io_axi_20_aw_bits_cache,io_axi_20_aw_bits_id,io_axi_20_aw_bits_len,io_axi_20_aw_bits_lock,io_axi_20_aw_bits_prot,io_axi_20_aw_bits_qos,io_axi_20_aw_bits_region,io_axi_20_aw_bits_size},
        io_axi_20_aw_valid,
        io_axi_20_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_20_ar(
        clock,
        reset,
        {io_axi_20_ar_bits_addr,io_axi_20_ar_bits_burst,io_axi_20_ar_bits_cache,io_axi_20_ar_bits_id,io_axi_20_ar_bits_len,io_axi_20_ar_bits_lock,io_axi_20_ar_bits_prot,io_axi_20_ar_bits_qos,io_axi_20_ar_bits_region,io_axi_20_ar_bits_size},
        io_axi_20_ar_valid,
        io_axi_20_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_20_w(
        clock,
        reset,
        {io_axi_20_w_bits_data,io_axi_20_w_bits_last,io_axi_20_w_bits_strb},
        io_axi_20_w_valid,
        io_axi_20_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_20_r(
        clock,
        reset,
        {io_axi_20_r_bits_data,io_axi_20_r_bits_last,io_axi_20_r_bits_resp,io_axi_20_r_bits_id},
        io_axi_20_r_valid,
        io_axi_20_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_20_b(
        clock,
        reset,
        {io_axi_20_b_bits_id,io_axi_20_b_bits_resp},
        io_axi_20_b_valid,
        io_axi_20_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_21_aw(
        clock,
        reset,
        {io_axi_21_aw_bits_addr,io_axi_21_aw_bits_burst,io_axi_21_aw_bits_cache,io_axi_21_aw_bits_id,io_axi_21_aw_bits_len,io_axi_21_aw_bits_lock,io_axi_21_aw_bits_prot,io_axi_21_aw_bits_qos,io_axi_21_aw_bits_region,io_axi_21_aw_bits_size},
        io_axi_21_aw_valid,
        io_axi_21_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_21_ar(
        clock,
        reset,
        {io_axi_21_ar_bits_addr,io_axi_21_ar_bits_burst,io_axi_21_ar_bits_cache,io_axi_21_ar_bits_id,io_axi_21_ar_bits_len,io_axi_21_ar_bits_lock,io_axi_21_ar_bits_prot,io_axi_21_ar_bits_qos,io_axi_21_ar_bits_region,io_axi_21_ar_bits_size},
        io_axi_21_ar_valid,
        io_axi_21_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_21_w(
        clock,
        reset,
        {io_axi_21_w_bits_data,io_axi_21_w_bits_last,io_axi_21_w_bits_strb},
        io_axi_21_w_valid,
        io_axi_21_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_21_r(
        clock,
        reset,
        {io_axi_21_r_bits_data,io_axi_21_r_bits_last,io_axi_21_r_bits_resp,io_axi_21_r_bits_id},
        io_axi_21_r_valid,
        io_axi_21_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_21_b(
        clock,
        reset,
        {io_axi_21_b_bits_id,io_axi_21_b_bits_resp},
        io_axi_21_b_valid,
        io_axi_21_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_22_aw(
        clock,
        reset,
        {io_axi_22_aw_bits_addr,io_axi_22_aw_bits_burst,io_axi_22_aw_bits_cache,io_axi_22_aw_bits_id,io_axi_22_aw_bits_len,io_axi_22_aw_bits_lock,io_axi_22_aw_bits_prot,io_axi_22_aw_bits_qos,io_axi_22_aw_bits_region,io_axi_22_aw_bits_size},
        io_axi_22_aw_valid,
        io_axi_22_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_22_ar(
        clock,
        reset,
        {io_axi_22_ar_bits_addr,io_axi_22_ar_bits_burst,io_axi_22_ar_bits_cache,io_axi_22_ar_bits_id,io_axi_22_ar_bits_len,io_axi_22_ar_bits_lock,io_axi_22_ar_bits_prot,io_axi_22_ar_bits_qos,io_axi_22_ar_bits_region,io_axi_22_ar_bits_size},
        io_axi_22_ar_valid,
        io_axi_22_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_22_w(
        clock,
        reset,
        {io_axi_22_w_bits_data,io_axi_22_w_bits_last,io_axi_22_w_bits_strb},
        io_axi_22_w_valid,
        io_axi_22_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_22_r(
        clock,
        reset,
        {io_axi_22_r_bits_data,io_axi_22_r_bits_last,io_axi_22_r_bits_resp,io_axi_22_r_bits_id},
        io_axi_22_r_valid,
        io_axi_22_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_22_b(
        clock,
        reset,
        {io_axi_22_b_bits_id,io_axi_22_b_bits_resp},
        io_axi_22_b_valid,
        io_axi_22_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_23_aw(
        clock,
        reset,
        {io_axi_23_aw_bits_addr,io_axi_23_aw_bits_burst,io_axi_23_aw_bits_cache,io_axi_23_aw_bits_id,io_axi_23_aw_bits_len,io_axi_23_aw_bits_lock,io_axi_23_aw_bits_prot,io_axi_23_aw_bits_qos,io_axi_23_aw_bits_region,io_axi_23_aw_bits_size},
        io_axi_23_aw_valid,
        io_axi_23_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_23_ar(
        clock,
        reset,
        {io_axi_23_ar_bits_addr,io_axi_23_ar_bits_burst,io_axi_23_ar_bits_cache,io_axi_23_ar_bits_id,io_axi_23_ar_bits_len,io_axi_23_ar_bits_lock,io_axi_23_ar_bits_prot,io_axi_23_ar_bits_qos,io_axi_23_ar_bits_region,io_axi_23_ar_bits_size},
        io_axi_23_ar_valid,
        io_axi_23_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_23_w(
        clock,
        reset,
        {io_axi_23_w_bits_data,io_axi_23_w_bits_last,io_axi_23_w_bits_strb},
        io_axi_23_w_valid,
        io_axi_23_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_23_r(
        clock,
        reset,
        {io_axi_23_r_bits_data,io_axi_23_r_bits_last,io_axi_23_r_bits_resp,io_axi_23_r_bits_id},
        io_axi_23_r_valid,
        io_axi_23_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_23_b(
        clock,
        reset,
        {io_axi_23_b_bits_id,io_axi_23_b_bits_resp},
        io_axi_23_b_valid,
        io_axi_23_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_24_aw(
        clock,
        reset,
        {io_axi_24_aw_bits_addr,io_axi_24_aw_bits_burst,io_axi_24_aw_bits_cache,io_axi_24_aw_bits_id,io_axi_24_aw_bits_len,io_axi_24_aw_bits_lock,io_axi_24_aw_bits_prot,io_axi_24_aw_bits_qos,io_axi_24_aw_bits_region,io_axi_24_aw_bits_size},
        io_axi_24_aw_valid,
        io_axi_24_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_24_ar(
        clock,
        reset,
        {io_axi_24_ar_bits_addr,io_axi_24_ar_bits_burst,io_axi_24_ar_bits_cache,io_axi_24_ar_bits_id,io_axi_24_ar_bits_len,io_axi_24_ar_bits_lock,io_axi_24_ar_bits_prot,io_axi_24_ar_bits_qos,io_axi_24_ar_bits_region,io_axi_24_ar_bits_size},
        io_axi_24_ar_valid,
        io_axi_24_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_24_w(
        clock,
        reset,
        {io_axi_24_w_bits_data,io_axi_24_w_bits_last,io_axi_24_w_bits_strb},
        io_axi_24_w_valid,
        io_axi_24_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_24_r(
        clock,
        reset,
        {io_axi_24_r_bits_data,io_axi_24_r_bits_last,io_axi_24_r_bits_resp,io_axi_24_r_bits_id},
        io_axi_24_r_valid,
        io_axi_24_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_24_b(
        clock,
        reset,
        {io_axi_24_b_bits_id,io_axi_24_b_bits_resp},
        io_axi_24_b_valid,
        io_axi_24_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_25_aw(
        clock,
        reset,
        {io_axi_25_aw_bits_addr,io_axi_25_aw_bits_burst,io_axi_25_aw_bits_cache,io_axi_25_aw_bits_id,io_axi_25_aw_bits_len,io_axi_25_aw_bits_lock,io_axi_25_aw_bits_prot,io_axi_25_aw_bits_qos,io_axi_25_aw_bits_region,io_axi_25_aw_bits_size},
        io_axi_25_aw_valid,
        io_axi_25_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_25_ar(
        clock,
        reset,
        {io_axi_25_ar_bits_addr,io_axi_25_ar_bits_burst,io_axi_25_ar_bits_cache,io_axi_25_ar_bits_id,io_axi_25_ar_bits_len,io_axi_25_ar_bits_lock,io_axi_25_ar_bits_prot,io_axi_25_ar_bits_qos,io_axi_25_ar_bits_region,io_axi_25_ar_bits_size},
        io_axi_25_ar_valid,
        io_axi_25_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_25_w(
        clock,
        reset,
        {io_axi_25_w_bits_data,io_axi_25_w_bits_last,io_axi_25_w_bits_strb},
        io_axi_25_w_valid,
        io_axi_25_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_25_r(
        clock,
        reset,
        {io_axi_25_r_bits_data,io_axi_25_r_bits_last,io_axi_25_r_bits_resp,io_axi_25_r_bits_id},
        io_axi_25_r_valid,
        io_axi_25_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_25_b(
        clock,
        reset,
        {io_axi_25_b_bits_id,io_axi_25_b_bits_resp},
        io_axi_25_b_valid,
        io_axi_25_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_26_aw(
        clock,
        reset,
        {io_axi_26_aw_bits_addr,io_axi_26_aw_bits_burst,io_axi_26_aw_bits_cache,io_axi_26_aw_bits_id,io_axi_26_aw_bits_len,io_axi_26_aw_bits_lock,io_axi_26_aw_bits_prot,io_axi_26_aw_bits_qos,io_axi_26_aw_bits_region,io_axi_26_aw_bits_size},
        io_axi_26_aw_valid,
        io_axi_26_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_26_ar(
        clock,
        reset,
        {io_axi_26_ar_bits_addr,io_axi_26_ar_bits_burst,io_axi_26_ar_bits_cache,io_axi_26_ar_bits_id,io_axi_26_ar_bits_len,io_axi_26_ar_bits_lock,io_axi_26_ar_bits_prot,io_axi_26_ar_bits_qos,io_axi_26_ar_bits_region,io_axi_26_ar_bits_size},
        io_axi_26_ar_valid,
        io_axi_26_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_26_w(
        clock,
        reset,
        {io_axi_26_w_bits_data,io_axi_26_w_bits_last,io_axi_26_w_bits_strb},
        io_axi_26_w_valid,
        io_axi_26_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_26_r(
        clock,
        reset,
        {io_axi_26_r_bits_data,io_axi_26_r_bits_last,io_axi_26_r_bits_resp,io_axi_26_r_bits_id},
        io_axi_26_r_valid,
        io_axi_26_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_26_b(
        clock,
        reset,
        {io_axi_26_b_bits_id,io_axi_26_b_bits_resp},
        io_axi_26_b_valid,
        io_axi_26_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_27_aw(
        clock,
        reset,
        {io_axi_27_aw_bits_addr,io_axi_27_aw_bits_burst,io_axi_27_aw_bits_cache,io_axi_27_aw_bits_id,io_axi_27_aw_bits_len,io_axi_27_aw_bits_lock,io_axi_27_aw_bits_prot,io_axi_27_aw_bits_qos,io_axi_27_aw_bits_region,io_axi_27_aw_bits_size},
        io_axi_27_aw_valid,
        io_axi_27_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_27_ar(
        clock,
        reset,
        {io_axi_27_ar_bits_addr,io_axi_27_ar_bits_burst,io_axi_27_ar_bits_cache,io_axi_27_ar_bits_id,io_axi_27_ar_bits_len,io_axi_27_ar_bits_lock,io_axi_27_ar_bits_prot,io_axi_27_ar_bits_qos,io_axi_27_ar_bits_region,io_axi_27_ar_bits_size},
        io_axi_27_ar_valid,
        io_axi_27_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_27_w(
        clock,
        reset,
        {io_axi_27_w_bits_data,io_axi_27_w_bits_last,io_axi_27_w_bits_strb},
        io_axi_27_w_valid,
        io_axi_27_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_27_r(
        clock,
        reset,
        {io_axi_27_r_bits_data,io_axi_27_r_bits_last,io_axi_27_r_bits_resp,io_axi_27_r_bits_id},
        io_axi_27_r_valid,
        io_axi_27_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_27_b(
        clock,
        reset,
        {io_axi_27_b_bits_id,io_axi_27_b_bits_resp},
        io_axi_27_b_valid,
        io_axi_27_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_28_aw(
        clock,
        reset,
        {io_axi_28_aw_bits_addr,io_axi_28_aw_bits_burst,io_axi_28_aw_bits_cache,io_axi_28_aw_bits_id,io_axi_28_aw_bits_len,io_axi_28_aw_bits_lock,io_axi_28_aw_bits_prot,io_axi_28_aw_bits_qos,io_axi_28_aw_bits_region,io_axi_28_aw_bits_size},
        io_axi_28_aw_valid,
        io_axi_28_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_28_ar(
        clock,
        reset,
        {io_axi_28_ar_bits_addr,io_axi_28_ar_bits_burst,io_axi_28_ar_bits_cache,io_axi_28_ar_bits_id,io_axi_28_ar_bits_len,io_axi_28_ar_bits_lock,io_axi_28_ar_bits_prot,io_axi_28_ar_bits_qos,io_axi_28_ar_bits_region,io_axi_28_ar_bits_size},
        io_axi_28_ar_valid,
        io_axi_28_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_28_w(
        clock,
        reset,
        {io_axi_28_w_bits_data,io_axi_28_w_bits_last,io_axi_28_w_bits_strb},
        io_axi_28_w_valid,
        io_axi_28_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_28_r(
        clock,
        reset,
        {io_axi_28_r_bits_data,io_axi_28_r_bits_last,io_axi_28_r_bits_resp,io_axi_28_r_bits_id},
        io_axi_28_r_valid,
        io_axi_28_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_28_b(
        clock,
        reset,
        {io_axi_28_b_bits_id,io_axi_28_b_bits_resp},
        io_axi_28_b_valid,
        io_axi_28_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_29_aw(
        clock,
        reset,
        {io_axi_29_aw_bits_addr,io_axi_29_aw_bits_burst,io_axi_29_aw_bits_cache,io_axi_29_aw_bits_id,io_axi_29_aw_bits_len,io_axi_29_aw_bits_lock,io_axi_29_aw_bits_prot,io_axi_29_aw_bits_qos,io_axi_29_aw_bits_region,io_axi_29_aw_bits_size},
        io_axi_29_aw_valid,
        io_axi_29_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_29_ar(
        clock,
        reset,
        {io_axi_29_ar_bits_addr,io_axi_29_ar_bits_burst,io_axi_29_ar_bits_cache,io_axi_29_ar_bits_id,io_axi_29_ar_bits_len,io_axi_29_ar_bits_lock,io_axi_29_ar_bits_prot,io_axi_29_ar_bits_qos,io_axi_29_ar_bits_region,io_axi_29_ar_bits_size},
        io_axi_29_ar_valid,
        io_axi_29_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_29_w(
        clock,
        reset,
        {io_axi_29_w_bits_data,io_axi_29_w_bits_last,io_axi_29_w_bits_strb},
        io_axi_29_w_valid,
        io_axi_29_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_29_r(
        clock,
        reset,
        {io_axi_29_r_bits_data,io_axi_29_r_bits_last,io_axi_29_r_bits_resp,io_axi_29_r_bits_id},
        io_axi_29_r_valid,
        io_axi_29_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_29_b(
        clock,
        reset,
        {io_axi_29_b_bits_id,io_axi_29_b_bits_resp},
        io_axi_29_b_valid,
        io_axi_29_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_30_aw(
        clock,
        reset,
        {io_axi_30_aw_bits_addr,io_axi_30_aw_bits_burst,io_axi_30_aw_bits_cache,io_axi_30_aw_bits_id,io_axi_30_aw_bits_len,io_axi_30_aw_bits_lock,io_axi_30_aw_bits_prot,io_axi_30_aw_bits_qos,io_axi_30_aw_bits_region,io_axi_30_aw_bits_size},
        io_axi_30_aw_valid,
        io_axi_30_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_30_ar(
        clock,
        reset,
        {io_axi_30_ar_bits_addr,io_axi_30_ar_bits_burst,io_axi_30_ar_bits_cache,io_axi_30_ar_bits_id,io_axi_30_ar_bits_len,io_axi_30_ar_bits_lock,io_axi_30_ar_bits_prot,io_axi_30_ar_bits_qos,io_axi_30_ar_bits_region,io_axi_30_ar_bits_size},
        io_axi_30_ar_valid,
        io_axi_30_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_30_w(
        clock,
        reset,
        {io_axi_30_w_bits_data,io_axi_30_w_bits_last,io_axi_30_w_bits_strb},
        io_axi_30_w_valid,
        io_axi_30_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_30_r(
        clock,
        reset,
        {io_axi_30_r_bits_data,io_axi_30_r_bits_last,io_axi_30_r_bits_resp,io_axi_30_r_bits_id},
        io_axi_30_r_valid,
        io_axi_30_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_30_b(
        clock,
        reset,
        {io_axi_30_b_bits_id,io_axi_30_b_bits_resp},
        io_axi_30_b_valid,
        io_axi_30_b_ready
);
// id, resp
// 6'h0, 2'h0

OUT#(64)out_io_axi_31_aw(
        clock,
        reset,
        {io_axi_31_aw_bits_addr,io_axi_31_aw_bits_burst,io_axi_31_aw_bits_cache,io_axi_31_aw_bits_id,io_axi_31_aw_bits_len,io_axi_31_aw_bits_lock,io_axi_31_aw_bits_prot,io_axi_31_aw_bits_qos,io_axi_31_aw_bits_region,io_axi_31_aw_bits_size},
        io_axi_31_aw_valid,
        io_axi_31_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(64)out_io_axi_31_ar(
        clock,
        reset,
        {io_axi_31_ar_bits_addr,io_axi_31_ar_bits_burst,io_axi_31_ar_bits_cache,io_axi_31_ar_bits_id,io_axi_31_ar_bits_len,io_axi_31_ar_bits_lock,io_axi_31_ar_bits_prot,io_axi_31_ar_bits_qos,io_axi_31_ar_bits_region,io_axi_31_ar_bits_size},
        io_axi_31_ar_valid,
        io_axi_31_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 33'h0, 2'h0, 4'h0, 6'h0, 4'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

OUT#(289)out_io_axi_31_w(
        clock,
        reset,
        {io_axi_31_w_bits_data,io_axi_31_w_bits_last,io_axi_31_w_bits_strb},
        io_axi_31_w_valid,
        io_axi_31_w_ready
);
// data, last, strb
// 256'h0, 1'h0, 32'h0

IN#(265)in_io_axi_31_r(
        clock,
        reset,
        {io_axi_31_r_bits_data,io_axi_31_r_bits_last,io_axi_31_r_bits_resp,io_axi_31_r_bits_id},
        io_axi_31_r_valid,
        io_axi_31_r_ready
);
// data, last, resp, id
// 256'h0, 1'h0, 2'h0, 6'h0

IN#(8)in_io_axi_31_b(
        clock,
        reset,
        {io_axi_31_b_bits_id,io_axi_31_b_bits_resp},
        io_axi_31_b_valid,
        io_axi_31_b_ready
);
// id, resp
// 6'h0, 2'h0


HBMCompress HBMCompress_inst(
        .*
);


initial begin
        reset <= 1;
        clock = 1;
        #1000;
        reset <= 0;
        #100;
		out_io_axi_0_aw.start();
		out_io_axi_0_w.start();
		out_io_axi_0_ar.start();
		
		out_io_axi_1_ar.start();
		out_io_axi_2_ar.start();
		out_io_axi_3_ar.start();
        #50;
		io_start <= 1;
		#13000;
		io_start_compress	<= 1;
		in_io_axi_0_r.write_many({256'h0, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_1_r.write_many({256'h1, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_2_r.write_many({256'h2, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_3_r.write_many({256'h3, 1'h0, 2'h0, 6'h0}, 2048);

		in_io_axi_0_r.write_many({256'h0, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_1_r.write_many({256'h1, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_2_r.write_many({256'h2, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_3_r.write_many({256'h3, 1'h0, 2'h0, 6'h0}, 2048);

		in_io_axi_0_r.write_many({256'h0, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_1_r.write_many({256'h1, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_2_r.write_many({256'h2, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_3_r.write_many({256'h3, 1'h0, 2'h0, 6'h0}, 2048);

		in_io_axi_0_r.write_many({256'h0, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_1_r.write_many({256'h1, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_2_r.write_many({256'h2, 1'h0, 2'h0, 6'h0}, 2048);
		in_io_axi_3_r.write_many({256'h3, 1'h0, 2'h0, 6'h0}, 2048);

		// #120_000;
		// io_start_compress	<= 0;
		// #10;
		// io_start_compress	<= 1;
		// in_io_axi_0_r.write_many({256'h0, 1'h0, 2'h0, 6'h0}, 2048);
		// in_io_axi_1_r.write_many({256'h1, 1'h0, 2'h0, 6'h0}, 2048);
		// in_io_axi_2_r.write_many({256'h2, 1'h0, 2'h0, 6'h0}, 2048);
		// in_io_axi_3_r.write_many({256'h3, 1'h0, 2'h0, 6'h0}, 2048);

end
always #5 clock=~clock;

endmodule